// Benchmark "multiplier_60917881_sat" written by ABC on Fri Nov 11 15:29:43 2022

module multiplier_60917881_sat ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] ,
    sat  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] ,
    \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ;
  output sat;
  wire new_n42_, new_n43_, new_n44_, new_n45_, new_n46_, new_n47_, new_n48_,
    new_n49_, new_n50_, new_n51_, new_n52_, new_n53_, new_n54_, new_n55_,
    new_n56_, new_n57_, new_n58_, new_n59_, new_n60_, new_n61_, new_n62_,
    new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_,
    new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_,
    new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_, new_n83_,
    new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_,
    new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_,
    new_n98_, new_n99_, new_n100_, new_n101_, new_n102_, new_n103_,
    new_n104_, new_n105_, new_n106_, new_n107_, new_n108_, new_n109_,
    new_n110_, new_n111_, new_n112_, new_n113_, new_n114_, new_n115_,
    new_n116_, new_n117_, new_n118_, new_n119_, new_n120_, new_n121_,
    new_n122_, new_n123_, new_n124_, new_n125_, new_n126_, new_n127_,
    new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_,
    new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_,
    new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_,
    new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_,
    new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_;
  assign sat = (~new_n42_ ^ (new_n447_ ^ ((~\a[2]  | (~new_n448_ & new_n484_) | (new_n448_ & ~new_n484_)) & (new_n339_ | (\a[2]  & (new_n448_ | ~new_n484_) & (~new_n448_ | new_n484_)) | (~\a[2]  & (new_n448_ ^ new_n484_)))))) & new_n450_ & (new_n339_ ^ (\a[2]  ^ (~new_n448_ ^ new_n484_)));
  assign new_n42_ = ~new_n336_ ^ (~new_n43_ ^ ((~\a[20]  | (~new_n269_ & new_n338_) | (new_n269_ & ~new_n338_)) & (new_n257_ | (\a[20]  & (new_n269_ | ~new_n338_) & (~new_n269_ | new_n338_)) | (~\a[20]  & (new_n269_ ^ new_n338_)))));
  assign new_n43_ = new_n335_ ^ ((~\a[14]  ^ \a[20] ) ^ (\a[5]  ^ ((new_n44_ & \a[8] ) | (~new_n278_ & (~new_n44_ | ~\a[8] ) & (new_n44_ | \a[8] )))));
  assign new_n44_ = ((\a[11]  & ((~new_n277_ & ~\a[14] ) | (new_n277_ & \a[14] ) | ((~new_n275_ | ~\a[14] ) & (new_n276_ | (new_n275_ & \a[14] ) | (~new_n275_ & ~\a[14] )))) & ((~new_n277_ ^ ~\a[14] ) | (new_n275_ & \a[14] ) | (~new_n276_ & (~new_n275_ | ~\a[14] ) & (new_n275_ | \a[14] )))) | (((\a[11]  & (new_n276_ | (new_n275_ & \a[14] ) | (~new_n275_ & ~\a[14] )) & (~new_n276_ | (new_n275_ ^ \a[14] ))) | (~new_n45_ & (~\a[11]  | (~new_n276_ & (~new_n275_ | ~\a[14] ) & (new_n275_ | \a[14] )) | (new_n276_ & (~new_n275_ ^ \a[14] ))) & (\a[11]  | (~new_n276_ ^ (new_n275_ ^ \a[14] ))))) & (~\a[11]  | ((new_n277_ | \a[14] ) & (~new_n277_ | ~\a[14] ) & ((new_n275_ & \a[14] ) | (~new_n276_ & (~new_n275_ | ~\a[14] ) & (new_n275_ | \a[14] )))) | ((new_n277_ ^ ~\a[14] ) & (~new_n275_ | ~\a[14] ) & (new_n276_ | (new_n275_ & \a[14] ) | (~new_n275_ & ~\a[14] )))) & (\a[11]  | ((~new_n277_ ^ ~\a[14] ) ^ ((new_n275_ & \a[14] ) | (~new_n276_ & (~new_n275_ | ~\a[14] ) & (new_n275_ | \a[14] ))))))) ^ (\a[11]  ^ ((~new_n256_ ^ ~\a[14] ) ^ ((new_n277_ & \a[14] ) | ((new_n277_ | \a[14] ) & (~new_n277_ | ~\a[14] ) & ((new_n275_ & \a[14] ) | (~new_n276_ & (~new_n275_ | ~\a[14] ) & (new_n275_ | \a[14] )))))));
  assign new_n45_ = (~new_n46_ | ~\a[11] ) & ((new_n46_ & \a[11] ) | (~new_n46_ & ~\a[11] ) | ((~\a[11]  | ((~new_n167_ | ~\a[14] ) & (new_n167_ | \a[14] ) & ((new_n212_ & \a[14] ) | ((~new_n212_ | ~\a[14] ) & (new_n212_ | \a[14] ) & ((new_n213_ & \a[14] ) | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] )))))) | ((~new_n167_ ^ \a[14] ) & (~new_n212_ | ~\a[14] ) & ((new_n212_ & \a[14] ) | (~new_n212_ & ~\a[14] ) | ((~new_n213_ | ~\a[14] ) & (new_n168_ | (new_n213_ & \a[14] ) | (~new_n213_ & ~\a[14] )))))) & (((~\a[11]  | ((~new_n212_ | ~\a[14] ) & (new_n212_ | \a[14] ) & ((new_n213_ & \a[14] ) | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] )))) | ((~new_n212_ ^ \a[14] ) & (~new_n213_ | ~\a[14] ) & (new_n168_ | (new_n213_ & \a[14] ) | (~new_n213_ & ~\a[14] )))) & (((~\a[11]  | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] )) | (new_n168_ & (~new_n213_ ^ \a[14] ))) & (new_n214_ | (\a[11]  & (new_n168_ | (new_n213_ & \a[14] ) | (~new_n213_ & ~\a[14] )) & (~new_n168_ | (new_n213_ ^ \a[14] ))) | (~\a[11]  & (new_n168_ ^ (new_n213_ ^ \a[14] ))))) | (\a[11]  & ((new_n212_ & \a[14] ) | (~new_n212_ & ~\a[14] ) | ((~new_n213_ | ~\a[14] ) & (new_n168_ | (new_n213_ & \a[14] ) | (~new_n213_ & ~\a[14] )))) & ((new_n212_ ^ \a[14] ) | (new_n213_ & \a[14] ) | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] )))) | (~\a[11]  & ((~new_n212_ ^ \a[14] ) ^ ((new_n213_ & \a[14] ) | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] ))))))) | (\a[11]  & ((new_n167_ & \a[14] ) | (~new_n167_ & ~\a[14] ) | ((~new_n212_ | ~\a[14] ) & ((new_n212_ & \a[14] ) | (~new_n212_ & ~\a[14] ) | ((~new_n213_ | ~\a[14] ) & (new_n168_ | (new_n213_ & \a[14] ) | (~new_n213_ & ~\a[14] )))))) & ((new_n167_ ^ \a[14] ) | (new_n212_ & \a[14] ) | ((~new_n212_ | ~\a[14] ) & (new_n212_ | \a[14] ) & ((new_n213_ & \a[14] ) | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] )))))) | (~\a[11]  & ((~new_n167_ ^ \a[14] ) ^ ((new_n212_ & \a[14] ) | ((~new_n212_ | ~\a[14] ) & (new_n212_ | \a[14] ) & ((new_n213_ & \a[14] ) | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] ))))))))));
  assign new_n46_ = ((new_n167_ & \a[14] ) | ((~new_n167_ | ~\a[14] ) & (new_n167_ | \a[14] ) & ((new_n212_ & \a[14] ) | ((new_n212_ | \a[14] ) & (~new_n212_ | ~\a[14] ) & ((new_n213_ & \a[14] ) | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] ))))))) ^ (\a[14]  ^ (~new_n47_ ^ new_n160_));
  assign new_n47_ = (~new_n48_ | ~\a[17] ) & (new_n122_ | (new_n48_ & \a[17] ) | (~new_n48_ & ~\a[17] ));
  assign new_n48_ = new_n117_ ^ (new_n49_ | new_n85_);
  assign new_n49_ = ~new_n81_ & (~new_n77_ | ((new_n83_ | new_n84_) & (new_n50_ | (~new_n83_ & ~new_n84_) | (new_n83_ & new_n84_)))) & (new_n77_ | (~new_n83_ & ~new_n84_) | (~new_n50_ & (new_n83_ | new_n84_) & (~new_n83_ | ~new_n84_)));
  assign new_n50_ = ~new_n51_ & ~new_n76_;
  assign new_n51_ = new_n72_ & (new_n52_ | (new_n71_ & (new_n56_ | (new_n70_ & (new_n59_ | (~new_n62_ & new_n69_))))));
  assign new_n52_ = (~\a[23]  ^ (new_n55_ & (~new_n53_ | ~new_n54_))) & ((\b[4]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] )) | (\b[3]  & \a[23]  & \a[24] ));
  assign new_n53_ = (\a[20]  | \a[21] ) & (~\a[20]  | ~\a[21] ) & (\a[22]  | \a[23] ) & (~\a[22]  | ~\a[23] );
  assign new_n54_ = ((\b[5]  & \b[6] ) | ((~\b[5]  | ~\b[6] ) & (\b[5]  | \b[6] ) & ((\b[4]  & \b[5] ) | (((\b[3]  & \b[4] ) | ((\b[3]  | \b[4] ) & (~\b[3]  | ~\b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))) & (~\b[4]  | ~\b[5] ) & (\b[4]  | \b[5] ))))) ^ (\b[6]  ^ \b[7] );
  assign new_n55_ = (~\b[5]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & (~\b[6]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[7]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] ));
  assign new_n56_ = (~\a[23]  ^ (new_n58_ & (~new_n53_ | ~new_n57_))) & ((\b[3]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] )) | (\b[2]  & \a[23]  & \a[24] ));
  assign new_n57_ = (\b[5]  ^ \b[6] ) ^ ((\b[4]  & \b[5] ) | (((\b[3]  & \b[4] ) | ((\b[3]  | \b[4] ) & (~\b[3]  | ~\b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))) & (~\b[4]  | ~\b[5] ) & (\b[4]  | \b[5] )));
  assign new_n58_ = (~\b[4]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & (~\b[5]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[6]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] ));
  assign new_n59_ = (~\a[23]  ^ (new_n61_ & (~new_n53_ | ~new_n60_))) & ((\b[2]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] )) | (\b[1]  & \a[23]  & \a[24] ));
  assign new_n60_ = ((\b[3]  & \b[4] ) | ((\b[3]  | \b[4] ) & (~\b[3]  | ~\b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))) ^ (\b[4]  ^ \b[5] );
  assign new_n61_ = (~\b[3]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & (~\b[4]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[5]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] ));
  assign new_n62_ = (new_n65_ | (\a[23]  ^ (new_n64_ & (~new_n53_ | ~new_n63_)))) & ((~new_n66_ & (new_n67_ | ~new_n68_)) | (~new_n65_ & (~\a[23]  ^ (new_n64_ & (~new_n53_ | ~new_n63_)))) | (new_n65_ & (~\a[23]  | ~new_n64_ | (new_n53_ & new_n63_)) & (\a[23]  | (new_n64_ & (~new_n53_ | ~new_n63_)))));
  assign new_n63_ = (~\b[3]  ^ ~\b[4] ) ^ ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] )));
  assign new_n64_ = (~\b[2]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & (~\b[3]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[4]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] ));
  assign new_n65_ = (~\b[1]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~\b[0]  | ~\a[23]  | ~\a[24] );
  assign new_n66_ = \b[0]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] ) & (~\b[0]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[1]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] )) & ((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\b[0]  ^ \b[1] )) & \a[23]  & (~\b[0]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~\b[0]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & ((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] )) & (~\b[1]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ));
  assign new_n67_ = \a[23]  ^ (((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & (~\b[3]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] )) & (~\b[2]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )));
  assign new_n68_ = (\b[0]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] )) ^ ((~\b[0]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[1]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] )) & ((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\b[0]  ^ \b[1] )) & \a[23]  & (~\b[0]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~\b[0]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & ((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] )) & (~\b[1]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )));
  assign new_n69_ = (~\a[23]  ^ (new_n61_ & (~new_n53_ | ~new_n60_))) ^ ((\b[2]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] )) | (\b[1]  & \a[23]  & \a[24] ));
  assign new_n70_ = (~\a[23]  ^ (new_n58_ & (~new_n53_ | ~new_n57_))) ^ ((\b[3]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] )) | (\b[2]  & \a[23]  & \a[24] ));
  assign new_n71_ = (~\a[23]  ^ (new_n55_ & (~new_n53_ | ~new_n54_))) ^ ((\b[4]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] )) | (\b[3]  & \a[23]  & \a[24] ));
  assign new_n72_ = ~new_n75_ ^ (~\a[23]  ^ (new_n74_ & (~new_n53_ | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n73_ & (~\b[7]  ^ \b[8] )))));
  assign new_n73_ = (~\b[6]  | ~\b[7] ) & (((~\b[5]  | ~\b[6] ) & ((\b[5]  & \b[6] ) | (~\b[5]  & ~\b[6] ) | ((~\b[4]  | ~\b[5] ) & (((~\b[3]  | ~\b[4] ) & ((~\b[3]  & ~\b[4] ) | (\b[3]  & \b[4] ) | ((~\b[2]  | ~\b[3] ) & ((~\b[2]  & ~\b[3] ) | (\b[2]  & \b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] ))))) | (\b[4]  & \b[5] ) | (~\b[4]  & ~\b[5] ))))) | (\b[6]  & \b[7] ) | (~\b[6]  & ~\b[7] ));
  assign new_n74_ = (~\b[6]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & (~\b[7]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[8]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] ));
  assign new_n75_ = (~\b[5]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~\b[4]  | ~\a[23]  | ~\a[24] );
  assign new_n76_ = ~new_n75_ & (~\a[23]  ^ (new_n74_ & (~new_n53_ | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n73_ & (~\b[7]  ^ \b[8] )))));
  assign new_n77_ = ~new_n80_ ^ (~new_n78_ ^ \a[23] );
  assign new_n78_ = new_n79_ & (~new_n53_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (\b[7]  | \b[8] ) & (~\b[7]  | ~\b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n73_ | (~\b[7]  & ~\b[8] ) | (\b[7]  & \b[8] ))))));
  assign new_n79_ = (~\b[8]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & (~\b[9]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[10]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] ));
  assign new_n80_ = (~\b[7]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~\b[6]  | ~\a[23]  | ~\a[24] );
  assign new_n81_ = \a[20]  ^ (((new_n82_ ^ \b[12] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[11]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] )) & (~\b[12]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )));
  assign new_n82_ = (~\b[11]  | ~\b[12] ) & ((\b[11]  & \b[12] ) | (~\b[11]  & ~\b[12] ) | ((~\b[10]  | ~\b[11] ) & ((\b[10]  & \b[11] ) | (~\b[10]  & ~\b[11] ) | ((~\b[9]  | ~\b[10] ) & ((~\b[9]  & ~\b[10] ) | (\b[9]  & \b[10] ) | ((~\b[8]  | ~\b[9] ) & ((~\b[8]  & ~\b[9] ) | (\b[8]  & \b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n73_ | (~\b[7]  & ~\b[8] ) | (\b[7]  & \b[8] ))))))))));
  assign new_n83_ = \a[23]  ^ (((~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n73_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[7]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[21]  ^ ~\a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[8]  | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[9]  | (~\a[22]  ^ ~\a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )));
  assign new_n84_ = (~\b[6]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~\b[5]  | ~\a[23]  | ~\a[24] );
  assign new_n85_ = new_n86_ & ((~new_n115_ & (new_n50_ | (new_n83_ & new_n84_) | (~new_n83_ & ~new_n84_)) & (~new_n50_ | (new_n83_ ^ new_n84_))) | ((new_n87_ | (~new_n91_ & new_n114_)) & (new_n115_ | (~new_n50_ & (~new_n83_ | ~new_n84_) & (new_n83_ | new_n84_)) | (new_n50_ & (~new_n83_ ^ new_n84_))) & (~new_n115_ | (~new_n50_ ^ (new_n83_ ^ new_n84_)))));
  assign new_n86_ = ~new_n81_ ^ (new_n77_ ^ ((~new_n83_ & ~new_n84_) | ((new_n51_ | new_n76_) & (new_n83_ | new_n84_) & (~new_n83_ | ~new_n84_))));
  assign new_n87_ = ~new_n88_ & new_n90_;
  assign new_n88_ = \a[20]  ^ ((~new_n89_ | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[9]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] )) & (~\b[10]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[11]  | (~\a[19]  ^ ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )));
  assign new_n89_ = (\b[10]  ^ \b[11] ) ^ ((\b[9]  & \b[10] ) | ((\b[9]  | \b[10] ) & (~\b[9]  | ~\b[10] ) & ((\b[8]  & \b[9] ) | ((\b[8]  | \b[9] ) & (~\b[8]  | ~\b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (\b[7]  | \b[8] ) & (~\b[7]  | ~\b[8] )))))));
  assign new_n90_ = new_n72_ ^ (new_n52_ | (new_n71_ & (new_n56_ | (new_n70_ & (new_n59_ | (~new_n62_ & new_n69_))))));
  assign new_n91_ = (~new_n92_ | new_n111_) & (((~new_n93_ | new_n113_) & ((~new_n94_ & (new_n96_ | ~new_n110_)) | (new_n93_ & ~new_n113_) | (~new_n93_ & new_n113_))) | (new_n92_ & ~new_n111_) | (~new_n92_ & new_n111_));
  assign new_n92_ = new_n71_ ^ (new_n56_ | (new_n70_ & (new_n59_ | (~new_n62_ & new_n69_))));
  assign new_n93_ = new_n70_ ^ (new_n59_ | (~new_n62_ & new_n69_));
  assign new_n94_ = ~new_n95_ & (new_n62_ | ~new_n69_) & (~new_n62_ | new_n69_);
  assign new_n95_ = \a[20]  ^ ((~\b[6]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] )) & (~\b[7]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[8]  | (~\a[19]  ^ ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & ((~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n73_ & (~\b[7]  ^ \b[8] ))));
  assign new_n96_ = (new_n97_ | ~new_n98_) & ((~new_n97_ & new_n98_) | (new_n97_ & ~new_n98_) | ((~new_n99_ | new_n100_) & (((new_n101_ | ~new_n109_) & (new_n102_ | (~new_n101_ & new_n109_) | (new_n101_ & ~new_n109_))) | (~new_n99_ & new_n100_) | (new_n99_ & ~new_n100_))));
  assign new_n97_ = \a[20]  ^ ((~new_n54_ | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[5]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] )) & (~\b[6]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[7]  | (~\a[19]  ^ ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )));
  assign new_n98_ = (new_n66_ | (~new_n67_ & new_n68_)) ^ (~new_n65_ ^ (~\a[23]  ^ (new_n64_ & (~new_n53_ | ~new_n63_))));
  assign new_n99_ = ~new_n67_ ^ new_n68_;
  assign new_n100_ = \a[20]  ^ ((~new_n57_ | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[4]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] )) & (~\b[5]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[6]  | (~\a[19]  ^ ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )));
  assign new_n101_ = \a[20]  ^ ((~new_n60_ | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[3]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] )) & (~\b[4]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[5]  | (~\a[19]  ^ ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )));
  assign new_n102_ = (~new_n105_ | (\a[20]  ^ (new_n104_ & (~new_n63_ | ~new_n103_)))) & ((~new_n106_ & (new_n107_ | ~new_n108_)) | (new_n105_ & (~\a[20]  ^ (new_n104_ & (~new_n63_ | ~new_n103_)))) | (~new_n105_ & (~\a[20]  | ~new_n104_ | (new_n63_ & new_n103_)) & (\a[20]  | (new_n104_ & (~new_n63_ | ~new_n103_)))));
  assign new_n103_ = (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ) & (\a[19]  | \a[20] ) & (~\a[19]  | ~\a[20] );
  assign new_n104_ = (~\b[3]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[4]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & (~\b[2]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ));
  assign new_n105_ = ((\b[0]  & (\a[20]  ^ ~\a[21] ) & (\a[21]  | \a[22] ) & (~\a[21]  | ~\a[22] )) | (\b[1]  & (\a[20]  | \a[21] ) & (~\a[20]  | ~\a[21] ) & (\a[22]  ^ ~\a[23] )) | ((\b[0]  ^ \b[1] ) & (\a[20]  | \a[21] ) & (~\a[20]  | ~\a[21] ) & (\a[22]  | \a[23] ) & (~\a[22]  | ~\a[23] ))) ^ (\a[23]  & \b[0]  & (\a[20]  | \a[21] ) & (~\a[20]  | ~\a[21] ));
  assign new_n106_ = \b[0]  & (\a[20]  | \a[21] ) & (~\a[20]  | ~\a[21] ) & (~\b[0]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[1]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\b[0]  ^ \b[1] )) & \a[20]  & (~\b[0]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & (~\b[1]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[0]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ));
  assign new_n107_ = \a[20]  ^ (((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & (~\b[2]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[1]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] )));
  assign new_n108_ = (\b[0]  & (\a[20]  | \a[21] ) & (~\a[20]  | ~\a[21] )) ^ ((~\b[0]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[1]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\b[0]  ^ \b[1] )) & \a[20]  & (~\b[0]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & (~\b[1]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[0]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] )));
  assign new_n109_ = ((~\b[0]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & (~\b[1]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[2]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] )) & ((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))) ^ (~\a[23]  | ((~\b[0]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[1]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] )) & ((~\b[0]  ^ \b[1] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] )) & \a[23]  & (~\b[0]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ))));
  assign new_n110_ = ~new_n95_ ^ (~new_n62_ ^ new_n69_);
  assign new_n111_ = \a[20]  ^ (new_n112_ & (~new_n103_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n73_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n112_ = (~\b[9]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[10]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & (~\b[8]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ));
  assign new_n113_ = \a[20]  ^ (((~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n73_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[7]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] )) & (~\b[8]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[9]  | (~\a[19]  ^ ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )));
  assign new_n114_ = ~new_n88_ ^ new_n90_;
  assign new_n115_ = \a[20]  ^ ((~new_n116_ | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[10]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] )) & (~\b[11]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[12]  | (~\a[19]  ^ ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )));
  assign new_n116_ = (\b[11]  ^ \b[12] ) ^ ((\b[10]  & \b[11] ) | ((~\b[10]  | ~\b[11] ) & (\b[10]  | \b[11] ) & ((\b[9]  & \b[10] ) | ((\b[9]  | \b[10] ) & (~\b[9]  | ~\b[10] ) & ((\b[8]  & \b[9] ) | ((\b[8]  | \b[9] ) & (~\b[8]  | ~\b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (\b[7]  | \b[8] ) & (~\b[7]  | ~\b[8] )))))))));
  assign new_n117_ = ~new_n121_ ^ (new_n118_ ^ ((~new_n120_ & ~new_n80_) | ((new_n120_ | new_n80_) & (~new_n120_ | ~new_n80_) & ((~new_n83_ & ~new_n84_) | ((~new_n83_ | ~new_n84_) & (new_n83_ | new_n84_) & (new_n51_ | new_n76_))))));
  assign new_n118_ = (new_n119_ ^ ~\a[23] ) ^ ((\b[8]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] )) | (\b[7]  & \a[23]  & \a[24] ));
  assign new_n119_ = (~\b[9]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[21]  ^ ~\a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[10]  | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[11]  | (~\a[22]  ^ ~\a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~new_n89_ | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ));
  assign new_n120_ = ~new_n78_ ^ ~\a[23] ;
  assign new_n121_ = \a[20]  ^ (~\b[12]  | (((~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] )) & (new_n82_ | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ))));
  assign new_n122_ = (~new_n124_ | ~\a[17] ) & ((new_n124_ & \a[17] ) | (~new_n124_ & ~\a[17] ) | ((~\a[17]  | (new_n123_ & (new_n87_ | (~new_n91_ & new_n114_))) | (~new_n123_ & ~new_n87_ & (new_n91_ | ~new_n114_))) & (((new_n159_ | (~new_n91_ & new_n114_) | (new_n91_ & ~new_n114_)) & (new_n125_ | (~new_n159_ & (new_n91_ | ~new_n114_) & (~new_n91_ | new_n114_)) | (new_n159_ & (new_n91_ ^ new_n114_)))) | (\a[17]  & (~new_n123_ | (~new_n87_ & (new_n91_ | ~new_n114_))) & (new_n123_ | new_n87_ | (~new_n91_ & new_n114_))) | (~\a[17]  & (~new_n123_ ^ (new_n87_ | (~new_n91_ & new_n114_)))))));
  assign new_n123_ = ~new_n115_ ^ (~new_n50_ ^ (~new_n83_ ^ ~new_n84_));
  assign new_n124_ = new_n86_ ^ ((~new_n115_ & (new_n50_ | (new_n83_ & new_n84_) | (~new_n83_ & ~new_n84_)) & (~new_n50_ | (new_n83_ ^ new_n84_))) | ((new_n87_ | (~new_n91_ & new_n114_)) & (new_n115_ | (~new_n50_ & (~new_n83_ | ~new_n84_) & (new_n83_ | new_n84_)) | (new_n50_ & (~new_n83_ ^ new_n84_))) & (~new_n115_ | (~new_n50_ ^ (new_n83_ ^ new_n84_)))));
  assign new_n125_ = ~new_n126_ & (~new_n158_ | (~new_n129_ & (~new_n157_ | (~new_n131_ & (new_n133_ | ~new_n156_)))));
  assign new_n126_ = ~new_n128_ & (~new_n127_ | ((~new_n93_ | new_n113_) & ((~new_n94_ & (new_n96_ | ~new_n110_)) | (new_n93_ & ~new_n113_) | (~new_n93_ & new_n113_)))) & (new_n127_ | (new_n93_ & ~new_n113_) | ((new_n94_ | (~new_n96_ & new_n110_)) & (~new_n93_ | new_n113_) & (new_n93_ | ~new_n113_)));
  assign new_n127_ = ~new_n111_ ^ (new_n71_ ^ (new_n56_ | (new_n70_ & (new_n59_ | (~new_n62_ & new_n69_)))));
  assign new_n128_ = \a[17]  ^ (((new_n82_ ^ \b[12] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[12]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[11]  | (~\a[15]  ^ ~\a[16] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n129_ = ~new_n130_ & ((new_n93_ & ~new_n113_) | (~new_n93_ & new_n113_) | (~new_n94_ & (new_n96_ | ~new_n110_))) & ((new_n93_ ^ ~new_n113_) | new_n94_ | (~new_n96_ & new_n110_));
  assign new_n130_ = \a[17]  ^ ((~new_n116_ | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[11]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[12]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[10]  | (~\a[15]  ^ ~\a[16] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n131_ = ~new_n132_ & (new_n96_ | ~new_n110_) & (~new_n96_ | new_n110_);
  assign new_n132_ = \a[17]  ^ ((~new_n89_ | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[10]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[11]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[9]  | (~\a[15]  ^ ~\a[16] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n133_ = (~new_n135_ | new_n153_) & ((new_n135_ & ~new_n153_) | (~new_n135_ & new_n153_) | (~new_n136_ & (~new_n152_ | ((new_n155_ | (new_n134_ & ~new_n102_) | (~new_n134_ & new_n102_)) & (new_n138_ | (~new_n155_ & (~new_n134_ | new_n102_) & (new_n134_ | ~new_n102_)) | (new_n155_ & (~new_n134_ ^ ~new_n102_)))))));
  assign new_n134_ = ~new_n101_ ^ new_n109_;
  assign new_n135_ = (~new_n97_ ^ new_n98_) ^ ((new_n99_ & ~new_n100_) | (((~new_n101_ & new_n109_) | (~new_n102_ & (new_n101_ | ~new_n109_) & (~new_n101_ | new_n109_))) & (new_n99_ | ~new_n100_) & (~new_n99_ | new_n100_)));
  assign new_n136_ = ~new_n137_ & ((~new_n99_ & new_n100_) | (new_n99_ & ~new_n100_) | ((new_n101_ | ~new_n109_) & (new_n102_ | (~new_n101_ & new_n109_) | (new_n101_ & ~new_n109_)))) & ((~new_n99_ ^ new_n100_) | (~new_n101_ & new_n109_) | (~new_n102_ & (new_n101_ | ~new_n109_) & (~new_n101_ | new_n109_)));
  assign new_n137_ = \a[17]  ^ (((~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n73_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[9]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[7]  | (~\a[15]  ^ ~\a[16] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n138_ = (new_n139_ | ~new_n140_) & ((~new_n139_ & new_n140_) | (new_n139_ & ~new_n140_) | ((~new_n141_ | new_n142_) & (((new_n143_ | ~new_n151_) & (new_n144_ | (~new_n143_ & new_n151_) | (new_n143_ & ~new_n151_))) | (~new_n141_ & new_n142_) | (new_n141_ & ~new_n142_))));
  assign new_n139_ = \a[17]  ^ ((~new_n54_ | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[6]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[7]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[5]  | (~\a[15]  ^ ~\a[16] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n140_ = (new_n106_ | (~new_n107_ & new_n108_)) ^ (new_n105_ ^ (~\a[20]  ^ (new_n104_ & (~new_n63_ | ~new_n103_))));
  assign new_n141_ = ~new_n107_ ^ new_n108_;
  assign new_n142_ = \a[17]  ^ ((~new_n57_ | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[5]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[6]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[4]  | (~\a[15]  ^ ~\a[16] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n143_ = \a[17]  ^ ((~new_n60_ | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[4]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[5]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[3]  | (~\a[15]  ^ ~\a[16] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n144_ = (~new_n147_ | (\a[17]  ^ (new_n146_ & (~new_n63_ | ~new_n145_)))) & ((~new_n148_ & (new_n149_ | ~new_n150_)) | (new_n147_ & (~\a[17]  ^ (new_n146_ & (~new_n63_ | ~new_n145_)))) | (~new_n147_ & (~\a[17]  | ~new_n146_ | (new_n63_ & new_n145_)) & (\a[17]  | (new_n146_ & (~new_n63_ | ~new_n145_)))));
  assign new_n145_ = (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ) & (\a[16]  | \a[17] ) & (~\a[16]  | ~\a[17] );
  assign new_n146_ = (~\b[3]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[4]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & (~\b[2]  | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ));
  assign new_n147_ = ((\b[0]  & (\a[17]  ^ ~\a[18] ) & (\a[18]  | \a[19] ) & (~\a[18]  | ~\a[19] )) | (\b[1]  & (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ) & (\a[19]  ^ ~\a[20] )) | ((\b[0]  ^ \b[1] ) & (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ) & (\a[19]  | \a[20] ) & (~\a[19]  | ~\a[20] ))) ^ (\a[20]  & \b[0]  & (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ));
  assign new_n148_ = \b[0]  & (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ) & (~\b[0]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[1]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\b[0]  ^ \b[1] )) & \a[17]  & (~\b[0]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & (~\b[1]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[0]  | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ));
  assign new_n149_ = \a[17]  ^ (((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & (~\b[2]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[1]  | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] )));
  assign new_n150_ = (\b[0]  & (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] )) ^ ((~\b[0]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[1]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\b[0]  ^ \b[1] )) & \a[17]  & (~\b[0]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & (~\b[1]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[0]  | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] )));
  assign new_n151_ = (~\a[20]  | ((~\b[0]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[1]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & ((~\b[0]  ^ \b[1] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] )) & \a[20]  & (~\b[0]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )))) ^ ((~\b[0]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] )) & (~\b[1]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[2]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n152_ = ~new_n137_ ^ ((~new_n99_ ^ new_n100_) ^ ((~new_n101_ & new_n109_) | (~new_n102_ & (new_n101_ | ~new_n109_) & (~new_n101_ | new_n109_))));
  assign new_n153_ = \a[17]  ^ (new_n154_ & (~new_n145_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n73_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n154_ = (~\b[9]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[10]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & (~\b[8]  | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ));
  assign new_n155_ = \a[17]  ^ (((~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n73_ & (~\b[7]  ^ \b[8] ))) & (~\b[7]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[8]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[6]  | (~\a[15]  ^ ~\a[16] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n156_ = ~new_n132_ ^ (~new_n96_ ^ new_n110_);
  assign new_n157_ = ~new_n130_ ^ ((new_n93_ ^ ~new_n113_) ^ (new_n94_ | (~new_n96_ & new_n110_)));
  assign new_n158_ = ~new_n128_ ^ (new_n127_ ^ ((new_n93_ & ~new_n113_) | ((new_n94_ | (~new_n96_ & new_n110_)) & (~new_n93_ | new_n113_) & (new_n93_ | ~new_n113_))));
  assign new_n159_ = \a[17]  ^ (~\b[12]  | ((new_n82_ | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & ((~\a[15]  ^ ~\a[16] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] ))));
  assign new_n160_ = \a[17]  ^ (new_n161_ ^ ((~new_n121_ & (new_n166_ | ~new_n118_) & (~new_n166_ | new_n118_)) | ((new_n49_ | new_n85_) & (new_n121_ | (~new_n166_ & new_n118_) | (new_n166_ & ~new_n118_)) & (~new_n121_ | (~new_n166_ ^ new_n118_)))));
  assign new_n161_ = \a[20]  ^ (~new_n162_ ^ new_n164_);
  assign new_n162_ = ~new_n163_ & (~new_n118_ | ((new_n120_ | new_n80_) & ((new_n120_ & new_n80_) | (~new_n120_ & ~new_n80_) | ((new_n83_ | new_n84_) & ((new_n83_ & new_n84_) | (~new_n83_ & ~new_n84_) | (~new_n51_ & ~new_n76_))))));
  assign new_n163_ = (new_n119_ ^ ~\a[23] ) & ((\b[8]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] )) | (\b[7]  & \a[23]  & \a[24] ));
  assign new_n164_ = (new_n165_ ^ ~\a[23] ) ^ ((\b[9]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] )) | (\b[8]  & \a[23]  & \a[24] ));
  assign new_n165_ = (~\b[10]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[21]  ^ ~\a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[11]  | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[12]  | (~\a[22]  ^ ~\a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~new_n116_ | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ));
  assign new_n166_ = (new_n120_ | new_n80_) & (~new_n77_ | ((new_n83_ | new_n84_) & (new_n50_ | (~new_n83_ & ~new_n84_) | (new_n83_ & new_n84_))));
  assign new_n167_ = ~new_n122_ ^ (new_n48_ ^ \a[17] );
  assign new_n168_ = (new_n171_ | ~new_n211_) & (~new_n169_ | ~\a[14] );
  assign new_n169_ = ~new_n125_ ^ new_n170_;
  assign new_n170_ = ~new_n159_ ^ (~new_n91_ ^ new_n114_);
  assign new_n171_ = (~new_n172_ | ~\a[14] ) & (((~new_n173_ | ~\a[14] ) & ((new_n173_ & \a[14] ) | (~new_n173_ & ~\a[14] ) | (~new_n174_ & (new_n176_ | new_n210_)))) | (new_n172_ & \a[14] ) | (~new_n172_ & ~\a[14] ));
  assign new_n172_ = new_n158_ ^ (new_n129_ | (new_n157_ & (new_n131_ | (~new_n133_ & new_n156_))));
  assign new_n173_ = new_n157_ ^ (new_n131_ | (~new_n133_ & new_n156_));
  assign new_n174_ = ~new_n175_ & (new_n133_ | ~new_n156_) & (~new_n133_ | new_n156_);
  assign new_n175_ = \a[14]  ^ (~\b[12]  | ((new_n82_ | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((~\a[12]  ^ ~\a[13] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  ^ ~\a[12] ))));
  assign new_n176_ = (~new_n177_ | new_n209_) & ((~new_n179_ & (~new_n208_ | (~new_n181_ & (new_n184_ | ~new_n207_)))) | (new_n177_ & ~new_n209_) | (~new_n177_ & new_n209_));
  assign new_n177_ = new_n178_ ^ (new_n136_ | (new_n152_ & ((~new_n155_ & (new_n102_ | (~new_n101_ & new_n109_) | (new_n101_ & ~new_n109_)) & (~new_n102_ | (~new_n101_ ^ new_n109_))) | (~new_n138_ & (new_n155_ | (~new_n102_ & (new_n101_ | ~new_n109_) & (~new_n101_ | new_n109_)) | (new_n102_ & (new_n101_ ^ new_n109_))) & (~new_n155_ | (~new_n102_ ^ (~new_n101_ ^ new_n109_)))))));
  assign new_n178_ = ~new_n153_ ^ ((~new_n97_ ^ new_n98_) ^ ((new_n99_ & ~new_n100_) | ((new_n99_ | ~new_n100_) & (~new_n99_ | new_n100_) & ((~new_n101_ & new_n109_) | (~new_n102_ & (new_n101_ | ~new_n109_) & (~new_n101_ | new_n109_))))));
  assign new_n179_ = ~new_n180_ & (~new_n152_ | ((new_n155_ | (~new_n102_ & (new_n101_ | ~new_n109_) & (~new_n101_ | new_n109_)) | (new_n102_ & (new_n101_ ^ new_n109_))) & (new_n138_ | (~new_n155_ & (new_n102_ | (~new_n101_ & new_n109_) | (new_n101_ & ~new_n109_)) & (~new_n102_ | (~new_n101_ ^ new_n109_))) | (new_n155_ & (new_n102_ ^ (~new_n101_ ^ new_n109_)))))) & (new_n152_ | (~new_n155_ & (new_n102_ | (~new_n101_ & new_n109_) | (new_n101_ & ~new_n109_)) & (~new_n102_ | (~new_n101_ ^ new_n109_))) | (~new_n138_ & (new_n155_ | (~new_n102_ & (new_n101_ | ~new_n109_) & (~new_n101_ | new_n109_)) | (new_n102_ & (new_n101_ ^ new_n109_))) & (~new_n155_ | (~new_n102_ ^ (~new_n101_ ^ new_n109_)))));
  assign new_n180_ = \a[14]  ^ ((~new_n116_ | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[11]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[12]  | (~\a[13]  ^ ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[10]  | (~\a[12]  ^ ~\a[13] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n181_ = ~new_n183_ & (new_n138_ | ~new_n182_) & (~new_n138_ | new_n182_);
  assign new_n182_ = ~new_n155_ ^ (~new_n102_ ^ (~new_n101_ ^ new_n109_));
  assign new_n183_ = \a[14]  ^ ((~new_n89_ | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[10]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[11]  | (~\a[13]  ^ ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[9]  | (~\a[12]  ^ ~\a[13] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n184_ = (~new_n186_ | new_n204_) & ((new_n186_ & ~new_n204_) | (~new_n186_ & new_n204_) | (~new_n187_ & (~new_n203_ | ((new_n206_ | (new_n185_ & ~new_n144_) | (~new_n185_ & new_n144_)) & (new_n189_ | (~new_n206_ & (~new_n185_ | new_n144_) & (new_n185_ | ~new_n144_)) | (new_n206_ & (~new_n185_ ^ ~new_n144_)))))));
  assign new_n185_ = ~new_n143_ ^ new_n151_;
  assign new_n186_ = (~new_n139_ ^ new_n140_) ^ ((new_n141_ & ~new_n142_) | (((~new_n143_ & new_n151_) | (~new_n144_ & (new_n143_ | ~new_n151_) & (~new_n143_ | new_n151_))) & (new_n141_ | ~new_n142_) & (~new_n141_ | new_n142_)));
  assign new_n187_ = ~new_n188_ & ((~new_n141_ & new_n142_) | (new_n141_ & ~new_n142_) | ((new_n143_ | ~new_n151_) & (new_n144_ | (~new_n143_ & new_n151_) | (new_n143_ & ~new_n151_)))) & ((~new_n141_ ^ new_n142_) | (~new_n143_ & new_n151_) | (~new_n144_ & (new_n143_ | ~new_n151_) & (~new_n143_ | new_n151_)));
  assign new_n188_ = \a[14]  ^ (((~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n73_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[9]  | (~\a[13]  ^ ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[7]  | (~\a[12]  ^ ~\a[13] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n189_ = (new_n190_ | ~new_n191_) & ((~new_n190_ & new_n191_) | (new_n190_ & ~new_n191_) | ((~new_n192_ | new_n193_) & (((new_n194_ | ~new_n202_) & (new_n195_ | (~new_n194_ & new_n202_) | (new_n194_ & ~new_n202_))) | (~new_n192_ & new_n193_) | (new_n192_ & ~new_n193_))));
  assign new_n190_ = \a[14]  ^ ((~new_n54_ | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[6]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[7]  | (~\a[13]  ^ ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[5]  | (~\a[12]  ^ ~\a[13] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n191_ = (new_n148_ | (~new_n149_ & new_n150_)) ^ (new_n147_ ^ (~\a[17]  ^ (new_n146_ & (~new_n63_ | ~new_n145_))));
  assign new_n192_ = ~new_n149_ ^ new_n150_;
  assign new_n193_ = \a[14]  ^ ((~new_n57_ | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[5]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[6]  | (~\a[13]  ^ ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[4]  | (~\a[12]  ^ ~\a[13] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n194_ = \a[14]  ^ ((~new_n60_ | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[4]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[5]  | (~\a[13]  ^ ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[3]  | (~\a[12]  ^ ~\a[13] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n195_ = (~new_n198_ | (\a[14]  ^ (new_n197_ & (~new_n63_ | ~new_n196_)))) & ((~new_n199_ & (new_n200_ | ~new_n201_)) | (new_n198_ & (~\a[14]  ^ (new_n197_ & (~new_n63_ | ~new_n196_)))) | (~new_n198_ & (~\a[14]  | ~new_n197_ | (new_n63_ & new_n196_)) & (\a[14]  | (new_n197_ & (~new_n63_ | ~new_n196_)))));
  assign new_n196_ = (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ) & (\a[13]  | \a[14] ) & (~\a[13]  | ~\a[14] );
  assign new_n197_ = (~\b[3]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[4]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & (~\b[2]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ));
  assign new_n198_ = ((\b[0]  & (\a[14]  ^ ~\a[15] ) & (\a[15]  | \a[16] ) & (~\a[15]  | ~\a[16] )) | (\b[1]  & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ) & (\a[16]  ^ ~\a[17] )) | ((\b[0]  ^ \b[1] ) & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ) & (\a[16]  | \a[17] ) & (~\a[16]  | ~\a[17] ))) ^ (\a[17]  & \b[0]  & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ));
  assign new_n199_ = \b[0]  & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ) & (~\b[0]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[1]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\b[0]  ^ \b[1] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & (~\b[1]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[0]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ));
  assign new_n200_ = \a[14]  ^ (((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & (~\b[2]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[1]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] )));
  assign new_n201_ = (\b[0]  & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] )) ^ ((~\b[0]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[1]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\b[0]  ^ \b[1] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & (~\b[1]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[0]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] )));
  assign new_n202_ = (~\a[17]  | ((~\b[0]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[1]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & ((~\b[0]  ^ \b[1] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] )) & \a[17]  & (~\b[0]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )))) ^ ((~\b[1]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[2]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] )));
  assign new_n203_ = ~new_n188_ ^ ((~new_n141_ ^ new_n142_) ^ ((~new_n143_ & new_n151_) | (~new_n144_ & (new_n143_ | ~new_n151_) & (~new_n143_ | new_n151_))));
  assign new_n204_ = \a[14]  ^ (new_n205_ & (~new_n196_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n73_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n205_ = (~\b[9]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[10]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & (~\b[8]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ));
  assign new_n206_ = \a[14]  ^ (((~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n73_ & (~\b[7]  ^ \b[8] ))) & (~\b[7]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[8]  | (~\a[13]  ^ ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[6]  | (~\a[12]  ^ ~\a[13] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n207_ = ~new_n183_ ^ (~new_n138_ ^ new_n182_);
  assign new_n208_ = ~new_n180_ ^ (new_n152_ ^ ((~new_n155_ & (new_n102_ | (~new_n101_ & new_n109_) | (new_n101_ & ~new_n109_)) & (~new_n102_ | (~new_n101_ ^ new_n109_))) | (~new_n138_ & (new_n155_ | (~new_n102_ & (new_n101_ | ~new_n109_) & (~new_n101_ | new_n109_)) | (new_n102_ & (new_n101_ ^ new_n109_))) & (~new_n155_ | (~new_n102_ ^ (~new_n101_ ^ new_n109_))))));
  assign new_n209_ = \a[14]  ^ (((new_n82_ ^ \b[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[12]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[11]  | (~\a[12]  ^ ~\a[13] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n210_ = new_n175_ & (new_n133_ ^ new_n156_);
  assign new_n211_ = \a[14]  ^ (~new_n125_ ^ new_n170_);
  assign new_n212_ = (new_n124_ ^ \a[17] ) ^ ((\a[17]  & (~new_n123_ | (~new_n87_ & (new_n91_ | ~new_n114_))) & (new_n123_ | new_n87_ | (~new_n91_ & new_n114_))) | (((~new_n159_ & (new_n91_ | ~new_n114_) & (~new_n91_ | new_n114_)) | (~new_n125_ & (new_n159_ | (~new_n91_ & new_n114_) | (new_n91_ & ~new_n114_)) & (~new_n159_ | (~new_n91_ ^ new_n114_)))) & (~\a[17]  | (new_n123_ & (new_n87_ | (~new_n91_ & new_n114_))) | (~new_n123_ & ~new_n87_ & (new_n91_ | ~new_n114_))) & (\a[17]  | (new_n123_ ^ (new_n87_ | (~new_n91_ & new_n114_))))));
  assign new_n213_ = ((~new_n159_ & (new_n91_ | ~new_n114_) & (~new_n91_ | new_n114_)) | (~new_n125_ & (new_n159_ | (~new_n91_ & new_n114_) | (new_n91_ & ~new_n114_)) & (~new_n159_ | (~new_n91_ ^ new_n114_)))) ^ (\a[17]  ^ (new_n123_ ^ (new_n87_ | (~new_n91_ & new_n114_))));
  assign new_n214_ = (~\a[11]  | (~new_n171_ & new_n211_) | (new_n171_ & ~new_n211_)) & ((\a[11]  & (new_n171_ | ~new_n211_) & (~new_n171_ | new_n211_)) | (~\a[11]  & (new_n171_ ^ new_n211_)) | ((~new_n215_ | ~\a[11] ) & ((new_n215_ & \a[11] ) | (~new_n215_ & ~\a[11] ) | ((~new_n216_ | ~\a[11] ) & (((new_n217_ | ~\a[11] ) & (new_n219_ | (~new_n217_ & \a[11] ) | (new_n217_ & ~\a[11] ))) | (new_n216_ & \a[11] ) | (~new_n216_ & ~\a[11] ))))));
  assign new_n215_ = ((new_n173_ & \a[14] ) | ((~new_n173_ | ~\a[14] ) & (new_n173_ | \a[14] ) & (new_n174_ | (~new_n176_ & ~new_n210_)))) ^ (new_n172_ ^ \a[14] );
  assign new_n216_ = (new_n173_ ^ \a[14] ) ^ (new_n174_ | (~new_n176_ & ~new_n210_));
  assign new_n217_ = ~new_n176_ ^ ~new_n218_;
  assign new_n218_ = ~new_n175_ ^ (~new_n133_ ^ new_n156_);
  assign new_n219_ = (~new_n220_ | ~\a[11] ) & (((~\a[11]  | (new_n208_ & (new_n181_ | (~new_n184_ & new_n207_))) | (~new_n208_ & ~new_n181_ & (new_n184_ | ~new_n207_))) & (((new_n255_ | (~new_n184_ & new_n207_) | (new_n184_ & ~new_n207_)) & (new_n221_ | (~new_n255_ & (new_n184_ | ~new_n207_) & (~new_n184_ | new_n207_)) | (new_n255_ & (new_n184_ ^ new_n207_)))) | (\a[11]  & (~new_n208_ | (~new_n181_ & (new_n184_ | ~new_n207_))) & (new_n208_ | new_n181_ | (~new_n184_ & new_n207_))) | (~\a[11]  & (~new_n208_ ^ (new_n181_ | (~new_n184_ & new_n207_)))))) | (new_n220_ & \a[11] ) | (~new_n220_ & ~\a[11] ));
  assign new_n220_ = (new_n179_ | (new_n208_ & (new_n181_ | (~new_n184_ & new_n207_)))) ^ (new_n177_ ^ ~new_n209_);
  assign new_n221_ = (~new_n222_ | new_n254_) & ((~new_n224_ & (~new_n253_ | (~new_n226_ & (new_n229_ | ~new_n252_)))) | (new_n222_ & ~new_n254_) | (~new_n222_ & new_n254_));
  assign new_n222_ = new_n223_ ^ (new_n187_ | (new_n203_ & ((~new_n206_ & (new_n144_ | (~new_n143_ & new_n151_) | (new_n143_ & ~new_n151_)) & (~new_n144_ | (~new_n143_ ^ new_n151_))) | (~new_n189_ & (new_n206_ | (~new_n144_ & (new_n143_ | ~new_n151_) & (~new_n143_ | new_n151_)) | (new_n144_ & (new_n143_ ^ new_n151_))) & (~new_n206_ | (~new_n144_ ^ (~new_n143_ ^ new_n151_)))))));
  assign new_n223_ = ~new_n204_ ^ ((~new_n139_ ^ new_n140_) ^ ((new_n141_ & ~new_n142_) | ((new_n141_ | ~new_n142_) & (~new_n141_ | new_n142_) & ((~new_n143_ & new_n151_) | (~new_n144_ & (new_n143_ | ~new_n151_) & (~new_n143_ | new_n151_))))));
  assign new_n224_ = ~new_n225_ & (~new_n203_ | ((new_n206_ | (~new_n144_ & (new_n143_ | ~new_n151_) & (~new_n143_ | new_n151_)) | (new_n144_ & (new_n143_ ^ new_n151_))) & (new_n189_ | (~new_n206_ & (new_n144_ | (~new_n143_ & new_n151_) | (new_n143_ & ~new_n151_)) & (~new_n144_ | (~new_n143_ ^ new_n151_))) | (new_n206_ & (new_n144_ ^ (~new_n143_ ^ new_n151_)))))) & (new_n203_ | (~new_n206_ & (new_n144_ | (~new_n143_ & new_n151_) | (new_n143_ & ~new_n151_)) & (~new_n144_ | (~new_n143_ ^ new_n151_))) | (~new_n189_ & (new_n206_ | (~new_n144_ & (new_n143_ | ~new_n151_) & (~new_n143_ | new_n151_)) | (new_n144_ & (new_n143_ ^ new_n151_))) & (~new_n206_ | (~new_n144_ ^ (~new_n143_ ^ new_n151_)))));
  assign new_n225_ = \a[11]  ^ ((~new_n116_ | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[11]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[12]  | (~\a[10]  ^ ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[10]  | (~\a[9]  ^ ~\a[10] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n226_ = ~new_n228_ & (new_n189_ | ~new_n227_) & (~new_n189_ | new_n227_);
  assign new_n227_ = ~new_n206_ ^ (~new_n144_ ^ (~new_n143_ ^ new_n151_));
  assign new_n228_ = \a[11]  ^ ((~new_n89_ | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[10]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[11]  | (~\a[10]  ^ ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[9]  | (~\a[9]  ^ ~\a[10] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n229_ = (~new_n231_ | new_n249_) & ((new_n231_ & ~new_n249_) | (~new_n231_ & new_n249_) | (~new_n232_ & (~new_n248_ | ((new_n251_ | (new_n230_ & ~new_n195_) | (~new_n230_ & new_n195_)) & (new_n234_ | (~new_n251_ & (~new_n230_ | new_n195_) & (new_n230_ | ~new_n195_)) | (new_n251_ & (~new_n230_ ^ ~new_n195_)))))));
  assign new_n230_ = ~new_n194_ ^ new_n202_;
  assign new_n231_ = (~new_n190_ ^ new_n191_) ^ ((new_n192_ & ~new_n193_) | (((~new_n194_ & new_n202_) | (~new_n195_ & (new_n194_ | ~new_n202_) & (~new_n194_ | new_n202_))) & (new_n192_ | ~new_n193_) & (~new_n192_ | new_n193_)));
  assign new_n232_ = ~new_n233_ & ((~new_n192_ & new_n193_) | (new_n192_ & ~new_n193_) | ((new_n194_ | ~new_n202_) & (new_n195_ | (~new_n194_ & new_n202_) | (new_n194_ & ~new_n202_)))) & ((~new_n192_ ^ new_n193_) | (~new_n194_ & new_n202_) | (~new_n195_ & (new_n194_ | ~new_n202_) & (~new_n194_ | new_n202_)));
  assign new_n233_ = \a[11]  ^ (((~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n73_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[9]  | (~\a[10]  ^ ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[7]  | (~\a[9]  ^ ~\a[10] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n234_ = (new_n235_ | ~new_n236_) & ((~new_n235_ & new_n236_) | (new_n235_ & ~new_n236_) | ((~new_n237_ | new_n238_) & (((new_n239_ | ~new_n247_) & (new_n240_ | (~new_n239_ & new_n247_) | (new_n239_ & ~new_n247_))) | (~new_n237_ & new_n238_) | (new_n237_ & ~new_n238_))));
  assign new_n235_ = \a[11]  ^ ((~new_n54_ | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[6]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[7]  | (~\a[10]  ^ ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[5]  | (~\a[9]  ^ ~\a[10] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n236_ = (new_n199_ | (~new_n200_ & new_n201_)) ^ (new_n198_ ^ (~\a[14]  ^ (new_n197_ & (~new_n63_ | ~new_n196_))));
  assign new_n237_ = ~new_n200_ ^ new_n201_;
  assign new_n238_ = \a[11]  ^ ((~new_n57_ | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[5]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[6]  | (~\a[10]  ^ ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[4]  | (~\a[9]  ^ ~\a[10] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n239_ = \a[11]  ^ ((~new_n60_ | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[4]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[5]  | (~\a[10]  ^ ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[3]  | (~\a[9]  ^ ~\a[10] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n240_ = (~new_n243_ | (\a[11]  ^ (new_n242_ & (~new_n63_ | ~new_n241_)))) & ((~new_n244_ & (new_n245_ | ~new_n246_)) | (new_n243_ & (~\a[11]  ^ (new_n242_ & (~new_n63_ | ~new_n241_)))) | (~new_n243_ & (~\a[11]  | ~new_n242_ | (new_n63_ & new_n241_)) & (\a[11]  | (new_n242_ & (~new_n63_ | ~new_n241_)))));
  assign new_n241_ = (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] );
  assign new_n242_ = (~\b[3]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[4]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[2]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ));
  assign new_n243_ = ((\b[0]  & (\a[11]  ^ ~\a[12] ) & (\a[12]  | \a[13] ) & (~\a[12]  | ~\a[13] )) | (\b[1]  & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ) & (\a[13]  ^ ~\a[14] )) | ((\b[0]  ^ \b[1] ) & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ) & (\a[13]  | \a[14] ) & (~\a[13]  | ~\a[14] ))) ^ (\a[14]  & \b[0]  & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ));
  assign new_n244_ = \b[0]  & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ) & (~\b[0]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\b[0]  ^ \b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[1]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[0]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ));
  assign new_n245_ = \a[11]  ^ (((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[2]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] )));
  assign new_n246_ = (\b[0]  & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] )) ^ ((~\b[0]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\b[0]  ^ \b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[1]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[0]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] )));
  assign new_n247_ = (~\a[14]  | ((~\b[0]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[1]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & ((~\b[0]  ^ \b[1] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )))) ^ ((~\b[1]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[2]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] )));
  assign new_n248_ = ~new_n233_ ^ ((~new_n192_ ^ new_n193_) ^ ((~new_n194_ & new_n202_) | (~new_n195_ & (new_n194_ | ~new_n202_) & (~new_n194_ | new_n202_))));
  assign new_n249_ = \a[11]  ^ (new_n250_ & (~new_n241_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n73_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n250_ = (~\b[9]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[10]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[8]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ));
  assign new_n251_ = \a[11]  ^ (((~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n73_ & (~\b[7]  ^ \b[8] ))) & (~\b[7]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[8]  | (~\a[10]  ^ ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[6]  | (~\a[9]  ^ ~\a[10] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n252_ = ~new_n228_ ^ (~new_n189_ ^ new_n227_);
  assign new_n253_ = ~new_n225_ ^ (new_n203_ ^ ((~new_n206_ & (new_n144_ | (~new_n143_ & new_n151_) | (new_n143_ & ~new_n151_)) & (~new_n144_ | (~new_n143_ ^ new_n151_))) | (~new_n189_ & (new_n206_ | (~new_n144_ & (new_n143_ | ~new_n151_) & (~new_n143_ | new_n151_)) | (new_n144_ & (new_n143_ ^ new_n151_))) & (~new_n206_ | (~new_n144_ ^ (~new_n143_ ^ new_n151_))))));
  assign new_n254_ = \a[11]  ^ (((new_n82_ ^ \b[12] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[12]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[11]  | (~\a[9]  ^ ~\a[10] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n255_ = \a[11]  ^ (~\b[12]  | ((new_n82_ | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((~\a[9]  ^ ~\a[10] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] ))));
  assign new_n256_ = ((new_n271_ & \a[17] ) | ((~new_n271_ | ~\a[17] ) & (new_n271_ | \a[17] ) & ((new_n273_ & \a[17] ) | ((new_n274_ | (~new_n47_ & new_n160_)) & (~new_n273_ | ~\a[17] ) & (new_n273_ | \a[17] ))))) ^ (\a[17]  ^ (~new_n257_ ^ new_n268_));
  assign new_n257_ = (~new_n265_ | ~\a[20] ) & (new_n258_ | (~new_n265_ & ~\a[20] ) | (new_n265_ & \a[20] ));
  assign new_n258_ = (~new_n259_ | ~\a[20] ) & ((new_n259_ & \a[20] ) | (~new_n259_ & ~\a[20] ) | ((~new_n264_ | ~\a[20] ) & ((new_n264_ & \a[20] ) | (~new_n264_ & ~\a[20] ) | ((new_n121_ | (~new_n166_ & new_n118_) | (new_n166_ & ~new_n118_)) & ((~new_n49_ & ~new_n85_) | (~new_n121_ & (new_n166_ | ~new_n118_) & (~new_n166_ | new_n118_)) | (new_n121_ & (new_n166_ ^ new_n118_)))))));
  assign new_n259_ = (~new_n260_ & ~new_n263_) ^ (new_n262_ | (~new_n162_ & new_n164_));
  assign new_n260_ = (new_n261_ ^ ~\a[23] ) & ((\b[10]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] )) | (\b[9]  & \a[23]  & \a[24] ));
  assign new_n261_ = ((new_n82_ ^ \b[12] ) | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~\b[12]  | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[11]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[21]  ^ ~\a[22] ) | (~\a[20]  ^ ~\a[21] ));
  assign new_n262_ = (new_n165_ ^ ~\a[23] ) & ((\b[9]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] )) | (\b[8]  & \a[23]  & \a[24] ));
  assign new_n263_ = (new_n261_ | \a[23] ) & (~new_n261_ | ~\a[23] ) & (~\b[10]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~\b[9]  | ~\a[23]  | ~\a[24] );
  assign new_n264_ = ~new_n162_ ^ new_n164_;
  assign new_n265_ = new_n266_ ^ (new_n260_ | (~new_n260_ & ~new_n263_ & (new_n262_ | (~new_n162_ & new_n164_))));
  assign new_n266_ = (~new_n267_ ^ \a[23] ) ^ ((~\b[11]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~\b[10]  | ~\a[23]  | ~\a[24] ));
  assign new_n267_ = \b[12]  & (((\a[22]  | \a[23] ) & (~\a[22]  | ~\a[23] ) & (\a[21]  ^ ~\a[22] ) & (\a[20]  ^ ~\a[21] )) | (~new_n82_ & (\a[22]  | \a[23] ) & (~\a[22]  | ~\a[23] ) & (\a[20]  | \a[21] ) & (~\a[20]  | ~\a[21] )));
  assign new_n268_ = \a[20]  ^ (~new_n269_ ^ (\a[23]  ? ((~\a[24]  | ~\b[11] ) & (~\b[12]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ))) : (\a[24]  & \b[12] )));
  assign new_n269_ = ((~new_n267_ ^ \a[23] ) | ((~\b[11]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~\b[10]  | ~\a[23]  | ~\a[24] ))) & (new_n270_ | ((new_n267_ ^ \a[23] ) & ((\b[11]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] )) | (\b[10]  & \a[23]  & \a[24] ))) | ((new_n267_ | ~\a[23] ) & (~new_n267_ | \a[23] ) & (~\b[11]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~\b[10]  | ~\a[23]  | ~\a[24] )));
  assign new_n270_ = ~new_n260_ & (new_n260_ | new_n263_ | (~new_n262_ & (new_n162_ | ~new_n164_)));
  assign new_n271_ = (~new_n265_ ^ \a[20] ) ^ ((~new_n259_ | ~\a[20] ) & ((new_n259_ & \a[20] ) | (~new_n259_ & ~\a[20] ) | ((~new_n264_ | ~\a[20] ) & ((new_n264_ & \a[20] ) | (~new_n264_ & ~\a[20] ) | ((new_n121_ | (~new_n166_ & new_n118_) | (new_n166_ & ~new_n118_)) & (new_n272_ | (~new_n121_ & (new_n166_ | ~new_n118_) & (~new_n166_ | new_n118_)) | (new_n121_ & (new_n166_ ^ new_n118_))))))));
  assign new_n272_ = ~new_n49_ & ~new_n85_;
  assign new_n273_ = (new_n259_ ^ \a[20] ) ^ ((new_n264_ & \a[20] ) | ((~new_n264_ | ~\a[20] ) & (new_n264_ | \a[20] ) & ((~new_n121_ & (new_n166_ | ~new_n118_) & (~new_n166_ | new_n118_)) | ((new_n49_ | new_n85_) & (new_n121_ | (~new_n166_ & new_n118_) | (new_n166_ & ~new_n118_)) & (~new_n121_ | (~new_n166_ ^ new_n118_))))));
  assign new_n274_ = \a[17]  & (~new_n161_ | ((new_n121_ | (~new_n166_ & new_n118_) | (new_n166_ & ~new_n118_)) & ((~new_n49_ & ~new_n85_) | (~new_n121_ & (new_n166_ | ~new_n118_) & (~new_n166_ | new_n118_)) | (new_n121_ & (new_n166_ ^ new_n118_))))) & (new_n161_ | (~new_n121_ & (new_n166_ | ~new_n118_) & (~new_n166_ | new_n118_)) | ((new_n49_ | new_n85_) & (new_n121_ | (~new_n166_ & new_n118_) | (new_n166_ & ~new_n118_)) & (~new_n121_ | (~new_n166_ ^ new_n118_))));
  assign new_n275_ = (new_n273_ ^ \a[17] ) ^ (new_n274_ | (~new_n47_ & new_n160_));
  assign new_n276_ = (~\a[14]  | (~new_n47_ & new_n160_) | (new_n47_ & ~new_n160_)) & (((~new_n167_ | ~\a[14] ) & ((new_n167_ & \a[14] ) | (~new_n167_ & ~\a[14] ) | ((~new_n212_ | ~\a[14] ) & ((~new_n212_ & ~\a[14] ) | (new_n212_ & \a[14] ) | ((~new_n213_ | ~\a[14] ) & (new_n168_ | (new_n213_ & \a[14] ) | (~new_n213_ & ~\a[14] ))))))) | (\a[14]  & (new_n47_ | ~new_n160_) & (~new_n47_ | new_n160_)) | (~\a[14]  & (new_n47_ ^ new_n160_)));
  assign new_n277_ = (new_n271_ ^ \a[17] ) ^ ((new_n273_ & \a[17] ) | ((new_n274_ | (~new_n47_ & new_n160_)) & (~new_n273_ | ~\a[17] ) & (new_n273_ | \a[17] )));
  assign new_n278_ = (~\a[8]  | (new_n281_ & (new_n279_ | (~new_n45_ & new_n280_))) | (~new_n281_ & ~new_n279_ & (new_n45_ | ~new_n280_))) & (((~\a[8]  | (~new_n45_ & new_n280_) | (new_n45_ & ~new_n280_)) & (((~new_n282_ | ~\a[8] ) & ((new_n282_ & \a[8] ) | (~new_n282_ & ~\a[8] ) | ((~new_n283_ | ~\a[8] ) & (new_n286_ | (new_n283_ & \a[8] ) | (~new_n283_ & ~\a[8] ))))) | (\a[8]  & (new_n45_ | ~new_n280_) & (~new_n45_ | new_n280_)) | (~\a[8]  & (new_n45_ ^ new_n280_)))) | (\a[8]  & (~new_n281_ | (~new_n279_ & (new_n45_ | ~new_n280_))) & (new_n281_ | new_n279_ | (~new_n45_ & new_n280_))) | (~\a[8]  & (~new_n281_ ^ (new_n279_ | (~new_n45_ & new_n280_)))));
  assign new_n279_ = \a[11]  & (new_n276_ | (new_n275_ & \a[14] ) | (~new_n275_ & ~\a[14] )) & (~new_n276_ | (new_n275_ ^ \a[14] ));
  assign new_n280_ = \a[11]  ^ (~new_n276_ ^ (new_n275_ ^ \a[14] ));
  assign new_n281_ = \a[11]  ^ (((new_n275_ & \a[14] ) | (~new_n276_ & (~new_n275_ | ~\a[14] ) & (new_n275_ | \a[14] ))) ^ (new_n277_ ^ \a[14] ));
  assign new_n282_ = (new_n46_ ^ \a[11] ) ^ ((\a[11]  & ((new_n167_ & \a[14] ) | (~new_n167_ & ~\a[14] ) | ((~new_n212_ | ~\a[14] ) & ((new_n212_ & \a[14] ) | (~new_n212_ & ~\a[14] ) | ((~new_n213_ | ~\a[14] ) & (new_n168_ | (new_n213_ & \a[14] ) | (~new_n213_ & ~\a[14] )))))) & ((new_n167_ ^ \a[14] ) | (new_n212_ & \a[14] ) | ((~new_n212_ | ~\a[14] ) & (new_n212_ | \a[14] ) & ((new_n213_ & \a[14] ) | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] )))))) | (((\a[11]  & ((new_n212_ & \a[14] ) | (~new_n212_ & ~\a[14] ) | ((~new_n213_ | ~\a[14] ) & (new_n168_ | (new_n213_ & \a[14] ) | (~new_n213_ & ~\a[14] )))) & ((new_n212_ ^ \a[14] ) | (new_n213_ & \a[14] ) | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] )))) | (((\a[11]  & (new_n168_ | (new_n213_ & \a[14] ) | (~new_n213_ & ~\a[14] )) & (~new_n168_ | (new_n213_ ^ \a[14] ))) | (~new_n214_ & (~\a[11]  | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] )) | (new_n168_ & (~new_n213_ ^ \a[14] ))) & (\a[11]  | (~new_n168_ ^ (new_n213_ ^ \a[14] ))))) & (~\a[11]  | ((~new_n212_ | ~\a[14] ) & (new_n212_ | \a[14] ) & ((new_n213_ & \a[14] ) | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] )))) | ((~new_n212_ ^ \a[14] ) & (~new_n213_ | ~\a[14] ) & (new_n168_ | (new_n213_ & \a[14] ) | (~new_n213_ & ~\a[14] )))) & (\a[11]  | ((new_n212_ ^ \a[14] ) ^ ((new_n213_ & \a[14] ) | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] ))))))) & (~\a[11]  | ((~new_n167_ | ~\a[14] ) & (new_n167_ | \a[14] ) & ((new_n212_ & \a[14] ) | ((~new_n212_ | ~\a[14] ) & (new_n212_ | \a[14] ) & ((new_n213_ & \a[14] ) | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] )))))) | ((~new_n167_ ^ \a[14] ) & (~new_n212_ | ~\a[14] ) & ((new_n212_ & \a[14] ) | (~new_n212_ & ~\a[14] ) | ((~new_n213_ | ~\a[14] ) & (new_n168_ | (new_n213_ & \a[14] ) | (~new_n213_ & ~\a[14] )))))) & (\a[11]  | ((new_n167_ ^ \a[14] ) ^ ((new_n212_ & \a[14] ) | ((~new_n212_ | ~\a[14] ) & (new_n212_ | \a[14] ) & ((new_n213_ & \a[14] ) | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] )))))))));
  assign new_n283_ = ((\a[11]  & ((new_n212_ & \a[14] ) | (~new_n212_ & ~\a[14] ) | ((~new_n213_ | ~\a[14] ) & (new_n168_ | (~new_n213_ & ~\a[14] ) | (new_n213_ & \a[14] )))) & ((new_n212_ ^ \a[14] ) | (new_n213_ & \a[14] ) | (~new_n168_ & (new_n213_ | \a[14] ) & (~new_n213_ | ~\a[14] )))) | (~new_n284_ & (~\a[11]  | ((~new_n212_ | ~\a[14] ) & (new_n212_ | \a[14] ) & ((new_n213_ & \a[14] ) | (~new_n168_ & (new_n213_ | \a[14] ) & (~new_n213_ | ~\a[14] )))) | ((~new_n212_ ^ \a[14] ) & (~new_n213_ | ~\a[14] ) & (new_n168_ | (~new_n213_ & ~\a[14] ) | (new_n213_ & \a[14] )))) & (\a[11]  | ((new_n212_ ^ \a[14] ) ^ ((new_n213_ & \a[14] ) | (~new_n168_ & (new_n213_ | \a[14] ) & (~new_n213_ | ~\a[14] ))))))) ^ (\a[11]  ^ ((~new_n167_ ^ ~\a[14] ) ^ ((new_n212_ & \a[14] ) | ((~new_n212_ | ~\a[14] ) & (new_n212_ | \a[14] ) & ((new_n213_ & \a[14] ) | (~new_n168_ & (new_n213_ | \a[14] ) & (~new_n213_ | ~\a[14] )))))));
  assign new_n284_ = (new_n214_ | ~new_n285_) & (~\a[11]  | (~new_n168_ & (new_n213_ | \a[14] ) & (~new_n213_ | ~\a[14] )) | (new_n168_ & (new_n213_ ^ ~\a[14] )));
  assign new_n285_ = \a[11]  ^ ((new_n213_ ^ \a[14] ) ^ ((new_n169_ & \a[14] ) | (~new_n171_ & (new_n169_ | \a[14] ) & (~new_n169_ | ~\a[14] ))));
  assign new_n286_ = (~\a[8]  | (~new_n284_ & new_n287_) | (new_n284_ & ~new_n287_)) & (new_n288_ | (\a[8]  & (new_n284_ | ~new_n287_) & (~new_n284_ | new_n287_)) | (~\a[8]  & (new_n284_ ^ new_n287_)));
  assign new_n287_ = \a[11]  ^ ((~new_n212_ ^ ~\a[14] ) ^ ((new_n213_ & \a[14] ) | (~new_n168_ & (~new_n213_ | ~\a[14] ) & (new_n213_ | \a[14] ))));
  assign new_n288_ = (~\a[8]  | (~new_n214_ & new_n285_) | (new_n214_ & ~new_n285_)) & ((\a[8]  & (new_n214_ | ~new_n285_) & (~new_n214_ | new_n285_)) | (~\a[8]  & (new_n214_ ^ new_n285_)) | ((~new_n289_ | ~\a[8] ) & ((new_n289_ & \a[8] ) | (~new_n289_ & ~\a[8] ) | ((~new_n290_ | ~\a[8] ) & ((new_n290_ & \a[8] ) | (~new_n290_ & ~\a[8] ) | ((~new_n291_ | ~\a[8] ) & (new_n292_ | (~new_n291_ & ~\a[8] ) | (new_n291_ & \a[8] ))))))));
  assign new_n289_ = (\a[11]  ^ (~new_n171_ ^ new_n211_)) ^ ((new_n215_ & \a[11] ) | ((~new_n215_ | ~\a[11] ) & (new_n215_ | \a[11] ) & ((new_n216_ & \a[11] ) | (((~new_n217_ & \a[11] ) | (~new_n219_ & (new_n217_ | ~\a[11] ) & (~new_n217_ | \a[11] ))) & (~new_n216_ | ~\a[11] ) & (new_n216_ | \a[11] )))));
  assign new_n290_ = (new_n215_ ^ \a[11] ) ^ ((new_n216_ & \a[11] ) | ((new_n216_ | \a[11] ) & (~new_n216_ | ~\a[11] ) & ((~new_n217_ & \a[11] ) | (~new_n219_ & (new_n217_ | ~\a[11] ) & (~new_n217_ | \a[11] )))));
  assign new_n291_ = (new_n216_ ^ \a[11] ) ^ ((~new_n217_ & \a[11] ) | (~new_n219_ & (new_n217_ | ~\a[11] ) & (~new_n217_ | \a[11] )));
  assign new_n292_ = (~\a[8]  | (~new_n219_ & new_n293_) | (new_n219_ & ~new_n293_)) & ((\a[8]  & (new_n219_ | ~new_n293_) & (~new_n219_ | new_n293_)) | (~\a[8]  & (new_n219_ ^ new_n293_)) | ((~new_n294_ | ~\a[8] ) & ((new_n294_ & \a[8] ) | (~new_n294_ & ~\a[8] ) | ((~new_n295_ | ~\a[8] ) & ((new_n295_ & \a[8] ) | (~new_n295_ & ~\a[8] ) | ((~new_n296_ | ~\a[8] ) & (new_n298_ | (~new_n296_ & ~\a[8] ) | (new_n296_ & \a[8] ))))))));
  assign new_n293_ = \a[11]  ^ (new_n176_ ^ ~new_n218_);
  assign new_n294_ = ((\a[11]  & (~new_n208_ | (~new_n181_ & (new_n184_ | ~new_n207_))) & (new_n208_ | new_n181_ | (~new_n184_ & new_n207_))) | (((~new_n255_ & (new_n184_ | ~new_n207_) & (~new_n184_ | new_n207_)) | (~new_n221_ & (new_n255_ | (~new_n184_ & new_n207_) | (new_n184_ & ~new_n207_)) & (~new_n255_ | (~new_n184_ ^ new_n207_)))) & (~\a[11]  | (new_n208_ & (new_n181_ | (~new_n184_ & new_n207_))) | (~new_n208_ & ~new_n181_ & (new_n184_ | ~new_n207_))) & (\a[11]  | (new_n208_ ^ (new_n181_ | (~new_n184_ & new_n207_)))))) ^ (new_n220_ ^ \a[11] );
  assign new_n295_ = ((~new_n255_ & (new_n184_ | ~new_n207_) & (~new_n184_ | new_n207_)) | (~new_n221_ & (new_n255_ | (~new_n184_ & new_n207_) | (new_n184_ & ~new_n207_)) & (~new_n255_ | (~new_n184_ ^ new_n207_)))) ^ (\a[11]  ^ (new_n208_ ^ (new_n181_ | (~new_n184_ & new_n207_))));
  assign new_n296_ = ~new_n221_ ^ new_n297_;
  assign new_n297_ = ~new_n255_ ^ (~new_n184_ ^ new_n207_);
  assign new_n298_ = (~new_n299_ | ~\a[8] ) & (((~\a[8]  | (new_n253_ & (new_n226_ | (~new_n229_ & new_n252_))) | (~new_n253_ & ~new_n226_ & (new_n229_ | ~new_n252_))) & (((new_n334_ | (~new_n229_ & new_n252_) | (new_n229_ & ~new_n252_)) & (new_n300_ | (~new_n334_ & (new_n229_ | ~new_n252_) & (~new_n229_ | new_n252_)) | (new_n334_ & (new_n229_ ^ new_n252_)))) | (\a[8]  & (~new_n253_ | (~new_n226_ & (new_n229_ | ~new_n252_))) & (new_n253_ | new_n226_ | (~new_n229_ & new_n252_))) | (~\a[8]  & (~new_n253_ ^ (new_n226_ | (~new_n229_ & new_n252_)))))) | (new_n299_ & \a[8] ) | (~new_n299_ & ~\a[8] ));
  assign new_n299_ = (new_n224_ | (new_n253_ & (new_n226_ | (~new_n229_ & new_n252_)))) ^ (new_n222_ ^ ~new_n254_);
  assign new_n300_ = (~new_n301_ | new_n333_) & ((~new_n303_ & (~new_n332_ | (~new_n305_ & (new_n308_ | ~new_n331_)))) | (new_n301_ & ~new_n333_) | (~new_n301_ & new_n333_));
  assign new_n301_ = new_n302_ ^ (new_n232_ | (new_n248_ & ((~new_n251_ & (new_n195_ | (~new_n194_ & new_n202_) | (new_n194_ & ~new_n202_)) & (~new_n195_ | (~new_n194_ ^ new_n202_))) | (~new_n234_ & (new_n251_ | (~new_n195_ & (new_n194_ | ~new_n202_) & (~new_n194_ | new_n202_)) | (new_n195_ & (new_n194_ ^ new_n202_))) & (~new_n251_ | (~new_n195_ ^ (~new_n194_ ^ new_n202_)))))));
  assign new_n302_ = ~new_n249_ ^ ((~new_n190_ ^ new_n191_) ^ ((new_n192_ & ~new_n193_) | ((new_n192_ | ~new_n193_) & (~new_n192_ | new_n193_) & ((~new_n194_ & new_n202_) | (~new_n195_ & (new_n194_ | ~new_n202_) & (~new_n194_ | new_n202_))))));
  assign new_n303_ = ~new_n304_ & (~new_n248_ | ((new_n251_ | (~new_n195_ & (new_n194_ | ~new_n202_) & (~new_n194_ | new_n202_)) | (new_n195_ & (new_n194_ ^ new_n202_))) & (new_n234_ | (~new_n251_ & (new_n195_ | (~new_n194_ & new_n202_) | (new_n194_ & ~new_n202_)) & (~new_n195_ | (~new_n194_ ^ new_n202_))) | (new_n251_ & (new_n195_ ^ (~new_n194_ ^ new_n202_)))))) & (new_n248_ | (~new_n251_ & (new_n195_ | (~new_n194_ & new_n202_) | (new_n194_ & ~new_n202_)) & (~new_n195_ | (~new_n194_ ^ new_n202_))) | (~new_n234_ & (new_n251_ | (~new_n195_ & (new_n194_ | ~new_n202_) & (~new_n194_ | new_n202_)) | (new_n195_ & (new_n194_ ^ new_n202_))) & (~new_n251_ | (~new_n195_ ^ (~new_n194_ ^ new_n202_)))));
  assign new_n304_ = \a[8]  ^ ((~new_n116_ | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[11]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[12]  | (~\a[7]  ^ ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[10]  | (~\a[6]  ^ ~\a[7] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n305_ = ~new_n307_ & (new_n234_ | ~new_n306_) & (~new_n234_ | new_n306_);
  assign new_n306_ = ~new_n251_ ^ (~new_n195_ ^ (~new_n194_ ^ new_n202_));
  assign new_n307_ = \a[8]  ^ ((~new_n89_ | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[10]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[11]  | (~\a[7]  ^ ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[9]  | (~\a[6]  ^ ~\a[7] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n308_ = (~new_n310_ | new_n328_) & ((new_n310_ & ~new_n328_) | (~new_n310_ & new_n328_) | (~new_n311_ & (~new_n327_ | ((new_n330_ | (new_n309_ & ~new_n240_) | (~new_n309_ & new_n240_)) & (new_n313_ | (~new_n330_ & (~new_n309_ | new_n240_) & (new_n309_ | ~new_n240_)) | (new_n330_ & (~new_n309_ ^ ~new_n240_)))))));
  assign new_n309_ = ~new_n239_ ^ new_n247_;
  assign new_n310_ = (~new_n235_ ^ new_n236_) ^ ((new_n237_ & ~new_n238_) | (((~new_n239_ & new_n247_) | (~new_n240_ & (new_n239_ | ~new_n247_) & (~new_n239_ | new_n247_))) & (new_n237_ | ~new_n238_) & (~new_n237_ | new_n238_)));
  assign new_n311_ = ~new_n312_ & ((~new_n237_ & new_n238_) | (new_n237_ & ~new_n238_) | ((new_n239_ | ~new_n247_) & (new_n240_ | (~new_n239_ & new_n247_) | (new_n239_ & ~new_n247_)))) & ((~new_n237_ ^ new_n238_) | (~new_n239_ & new_n247_) | (~new_n240_ & (new_n239_ | ~new_n247_) & (~new_n239_ | new_n247_)));
  assign new_n312_ = \a[8]  ^ (((~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n73_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[9]  | (~\a[7]  ^ ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[7]  | (~\a[6]  ^ ~\a[7] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n313_ = (~new_n314_ | new_n315_) & ((~new_n314_ & new_n315_) | (new_n314_ & ~new_n315_) | ((~new_n316_ | new_n317_) & (((new_n318_ | ~new_n326_) & (new_n319_ | (~new_n318_ & new_n326_) | (new_n318_ & ~new_n326_))) | (~new_n316_ & new_n317_) | (new_n316_ & ~new_n317_))));
  assign new_n314_ = (new_n244_ | (~new_n245_ & new_n246_)) ^ (new_n243_ ^ (~\a[11]  ^ (new_n242_ & (~new_n63_ | ~new_n241_))));
  assign new_n315_ = \a[8]  ^ ((~new_n54_ | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[6]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[7]  | (~\a[7]  ^ ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[5]  | (~\a[6]  ^ ~\a[7] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n316_ = ~new_n245_ ^ new_n246_;
  assign new_n317_ = \a[8]  ^ ((~new_n57_ | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[5]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[6]  | (~\a[7]  ^ ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[4]  | (~\a[6]  ^ ~\a[7] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n318_ = \a[8]  ^ ((~new_n60_ | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[4]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[5]  | (~\a[7]  ^ ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[3]  | (~\a[6]  ^ ~\a[7] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n319_ = (~new_n322_ | (\a[8]  ^ (new_n321_ & (~new_n63_ | ~new_n320_)))) & ((~new_n323_ & (new_n324_ | ~new_n325_)) | (new_n322_ & (~\a[8]  ^ (new_n321_ & (~new_n63_ | ~new_n320_)))) | (~new_n322_ & (~\a[8]  | ~new_n321_ | (new_n63_ & new_n320_)) & (\a[8]  | (new_n321_ & (~new_n63_ | ~new_n320_)))));
  assign new_n320_ = (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] );
  assign new_n321_ = (~\b[3]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[4]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[2]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ));
  assign new_n322_ = ((\b[0]  & (\a[8]  ^ ~\a[9] ) & (\a[9]  | \a[10] ) & (~\a[9]  | ~\a[10] )) | (\b[1]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  ^ ~\a[11] )) | ((\b[0]  ^ \b[1] ) & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] ))) ^ (\a[11]  & \b[0]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ));
  assign new_n323_ = \b[0]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (~\b[0]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\b[0]  ^ \b[1] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[1]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ));
  assign new_n324_ = \a[8]  ^ (((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[2]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )));
  assign new_n325_ = (\b[0]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] )) ^ ((~\b[0]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\b[0]  ^ \b[1] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[1]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )));
  assign new_n326_ = (~\a[11]  | ((~\b[0]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\b[0]  ^ \b[1] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )))) ^ ((~\b[1]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[2]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] )));
  assign new_n327_ = ~new_n312_ ^ ((~new_n237_ ^ new_n238_) ^ ((~new_n239_ & new_n247_) | (~new_n240_ & (new_n239_ | ~new_n247_) & (~new_n239_ | new_n247_))));
  assign new_n328_ = \a[8]  ^ (new_n329_ & (~new_n320_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n73_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n329_ = (~\b[9]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[10]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[8]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ));
  assign new_n330_ = \a[8]  ^ (((~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n73_ & (~\b[7]  ^ \b[8] ))) & (~\b[7]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[8]  | (~\a[7]  ^ ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[6]  | (~\a[6]  ^ ~\a[7] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n331_ = ~new_n307_ ^ (~new_n234_ ^ new_n306_);
  assign new_n332_ = ~new_n304_ ^ (new_n248_ ^ ((~new_n251_ & (new_n195_ | (~new_n194_ & new_n202_) | (new_n194_ & ~new_n202_)) & (~new_n195_ | (~new_n194_ ^ new_n202_))) | (~new_n234_ & (new_n251_ | (~new_n195_ & (new_n194_ | ~new_n202_) & (~new_n194_ | new_n202_)) | (new_n195_ & (new_n194_ ^ new_n202_))) & (~new_n251_ | (~new_n195_ ^ (~new_n194_ ^ new_n202_))))));
  assign new_n333_ = \a[8]  ^ (((new_n82_ ^ \b[12] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[12]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[11]  | (~\a[6]  ^ ~\a[7] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n334_ = \a[8]  ^ (~\b[12]  | ((new_n82_ | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[6]  ^ ~\a[7] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  ^ ~\a[6] ))));
  assign new_n335_ = (~\a[17]  | (~new_n257_ & new_n268_) | (new_n257_ & ~new_n268_)) & (((~new_n271_ | ~\a[17] ) & ((new_n271_ & \a[17] ) | (~new_n271_ & ~\a[17] ) | ((~new_n273_ | ~\a[17] ) & ((~new_n274_ & (new_n47_ | ~new_n160_)) | (new_n273_ & \a[17] ) | (~new_n273_ & ~\a[17] ))))) | (\a[17]  & (new_n257_ | ~new_n268_) & (~new_n257_ | new_n268_)) | (~\a[17]  & (new_n257_ ^ new_n268_)));
  assign new_n336_ = ~new_n337_ ^ ((\a[23]  & (~\a[24]  | ~\b[12] )) ^ (\a[2]  ^ ((\a[23]  & ((\b[12]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] )) | (\a[24]  & \b[11] ))) | (~new_n269_ & (~\a[23]  | ((~\b[12]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~\a[24]  | ~\b[11] ))) & (\a[23]  | (\a[24]  & \b[12] ))))));
  assign new_n337_ = \a[17]  ^ ((\a[11]  & ((~new_n256_ & ~\a[14] ) | (new_n256_ & \a[14] ) | ((~new_n277_ | ~\a[14] ) & ((~new_n277_ & ~\a[14] ) | (new_n277_ & \a[14] ) | ((~new_n275_ | ~\a[14] ) & (new_n276_ | (new_n275_ & \a[14] ) | (~new_n275_ & ~\a[14] )))))) & ((~new_n256_ ^ ~\a[14] ) | (new_n277_ & \a[14] ) | ((new_n277_ | \a[14] ) & (~new_n277_ | ~\a[14] ) & ((new_n275_ & \a[14] ) | (~new_n276_ & (~new_n275_ | ~\a[14] ) & (new_n275_ | \a[14] )))))) | (((\a[11]  & ((~new_n277_ & ~\a[14] ) | (new_n277_ & \a[14] ) | ((~new_n275_ | ~\a[14] ) & (new_n276_ | (new_n275_ & \a[14] ) | (~new_n275_ & ~\a[14] )))) & ((~new_n277_ ^ ~\a[14] ) | (new_n275_ & \a[14] ) | (~new_n276_ & (~new_n275_ | ~\a[14] ) & (new_n275_ | \a[14] )))) | (((\a[11]  & (new_n276_ | (new_n275_ & \a[14] ) | (~new_n275_ & ~\a[14] )) & (~new_n276_ | (new_n275_ ^ \a[14] ))) | (~new_n45_ & (~\a[11]  | (~new_n276_ & (~new_n275_ | ~\a[14] ) & (new_n275_ | \a[14] )) | (new_n276_ & (~new_n275_ ^ \a[14] ))) & (\a[11]  | (~new_n276_ ^ (new_n275_ ^ \a[14] ))))) & (~\a[11]  | ((new_n277_ | \a[14] ) & (~new_n277_ | ~\a[14] ) & ((new_n275_ & \a[14] ) | (~new_n276_ & (~new_n275_ | ~\a[14] ) & (new_n275_ | \a[14] )))) | ((new_n277_ ^ ~\a[14] ) & (~new_n275_ | ~\a[14] ) & (new_n276_ | (new_n275_ & \a[14] ) | (~new_n275_ & ~\a[14] )))) & (\a[11]  | ((~new_n277_ ^ ~\a[14] ) ^ ((new_n275_ & \a[14] ) | (~new_n276_ & (~new_n275_ | ~\a[14] ) & (new_n275_ | \a[14] ))))))) & (~\a[11]  | ((new_n256_ | \a[14] ) & (~new_n256_ | ~\a[14] ) & ((new_n277_ & \a[14] ) | ((new_n277_ | \a[14] ) & (~new_n277_ | ~\a[14] ) & ((new_n275_ & \a[14] ) | (~new_n276_ & (~new_n275_ | ~\a[14] ) & (new_n275_ | \a[14] )))))) | ((new_n256_ ^ ~\a[14] ) & (~new_n277_ | ~\a[14] ) & ((~new_n277_ & ~\a[14] ) | (new_n277_ & \a[14] ) | ((~new_n275_ | ~\a[14] ) & (new_n276_ | (new_n275_ & \a[14] ) | (~new_n275_ & ~\a[14] )))))) & (\a[11]  | ((~new_n256_ ^ ~\a[14] ) ^ ((new_n277_ & \a[14] ) | ((new_n277_ | \a[14] ) & (~new_n277_ | ~\a[14] ) & ((new_n275_ & \a[14] ) | (~new_n276_ & (~new_n275_ | ~\a[14] ) & (new_n275_ | \a[14] )))))))));
  assign new_n338_ = \a[23]  ? ((~\a[24]  | ~\b[11] ) & (~\b[12]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ))) : (\a[24]  & \b[12] );
  assign new_n339_ = (~new_n340_ | ~\a[2] ) & ((new_n340_ & \a[2] ) | (~new_n340_ & ~\a[2] ) | ((~new_n393_ | ~\a[2] ) & ((~new_n393_ & ~\a[2] ) | (new_n393_ & \a[2] ) | ((~new_n394_ | ~\a[2] ) & ((new_n394_ & \a[2] ) | (~new_n394_ & ~\a[2] ) | ((~\a[2]  | (~new_n345_ & new_n392_) | (new_n345_ & ~new_n392_)) & (new_n395_ | (\a[2]  & (new_n345_ | ~new_n392_) & (~new_n345_ | new_n392_)) | (~\a[2]  & (new_n345_ ^ new_n392_)))))))));
  assign new_n340_ = (new_n341_ ^ \a[5] ) ^ ((new_n342_ & \a[5] ) | ((new_n342_ | \a[5] ) & (~new_n342_ | ~\a[5] ) & ((new_n343_ & \a[5] ) | ((~new_n343_ | ~\a[5] ) & (new_n343_ | \a[5] ) & (new_n344_ | (~new_n345_ & new_n392_))))));
  assign new_n341_ = ((\a[8]  & (new_n45_ | ~new_n280_) & (~new_n45_ | new_n280_)) | (((new_n282_ & \a[8] ) | ((~new_n282_ | ~\a[8] ) & (new_n282_ | \a[8] ) & ((new_n283_ & \a[8] ) | (~new_n286_ & (~new_n283_ | ~\a[8] ) & (new_n283_ | \a[8] ))))) & (~\a[8]  | (~new_n45_ & new_n280_) | (new_n45_ & ~new_n280_)) & (\a[8]  | (~new_n45_ ^ new_n280_)))) ^ (\a[8]  ^ (new_n281_ ^ (new_n279_ | (~new_n45_ & new_n280_))));
  assign new_n342_ = ((new_n282_ & \a[8] ) | (((new_n283_ & \a[8] ) | (~new_n286_ & (new_n283_ | \a[8] ) & (~new_n283_ | ~\a[8] ))) & (new_n282_ | \a[8] ) & (~new_n282_ | ~\a[8] ))) ^ (\a[8]  ^ (~new_n45_ ^ new_n280_));
  assign new_n343_ = (new_n282_ ^ \a[8] ) ^ ((new_n283_ & \a[8] ) | (~new_n286_ & (~new_n283_ | ~\a[8] ) & (new_n283_ | \a[8] )));
  assign new_n344_ = \a[5]  & (new_n286_ | (new_n283_ & \a[8] ) | (~new_n283_ & ~\a[8] )) & (~new_n286_ | (new_n283_ ^ \a[8] ));
  assign new_n345_ = (~new_n346_ | ~\a[5] ) & (new_n347_ | (new_n346_ & \a[5] ) | (~new_n346_ & ~\a[5] ));
  assign new_n346_ = ~new_n288_ ^ (\a[8]  ^ (~new_n284_ ^ new_n287_));
  assign new_n347_ = (~\a[5]  | ((~new_n348_ | ~\a[8] ) & (new_n348_ | \a[8] ) & ((new_n289_ & \a[8] ) | ((~new_n289_ | ~\a[8] ) & (new_n289_ | \a[8] ) & ((new_n290_ & \a[8] ) | ((~new_n290_ | ~\a[8] ) & (new_n290_ | \a[8] ) & ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))))))) | ((~new_n348_ ^ \a[8] ) & (~new_n289_ | ~\a[8] ) & ((new_n289_ & \a[8] ) | (~new_n289_ & ~\a[8] ) | ((~new_n290_ | ~\a[8] ) & ((new_n290_ & \a[8] ) | (~new_n290_ & ~\a[8] ) | ((~new_n291_ | ~\a[8] ) & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )))))))) & (((~\a[5]  | ((~new_n289_ | ~\a[8] ) & (new_n289_ | \a[8] ) & ((new_n290_ & \a[8] ) | ((~new_n290_ | ~\a[8] ) & (new_n290_ | \a[8] ) & ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))))) | ((~new_n289_ ^ \a[8] ) & (~new_n290_ | ~\a[8] ) & ((new_n290_ & \a[8] ) | (~new_n290_ & ~\a[8] ) | ((~new_n291_ | ~\a[8] ) & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )))))) & ((\a[5]  & ((new_n289_ & \a[8] ) | (~new_n289_ & ~\a[8] ) | ((~new_n290_ | ~\a[8] ) & ((new_n290_ & \a[8] ) | (~new_n290_ & ~\a[8] ) | ((~new_n291_ | ~\a[8] ) & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )))))) & ((new_n289_ ^ \a[8] ) | (new_n290_ & \a[8] ) | ((~new_n290_ | ~\a[8] ) & (new_n290_ | \a[8] ) & ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))))) | (~\a[5]  & ((~new_n289_ ^ \a[8] ) ^ ((new_n290_ & \a[8] ) | ((~new_n290_ | ~\a[8] ) & (new_n290_ | \a[8] ) & ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] ))))))) | ((~\a[5]  | ((~new_n290_ | ~\a[8] ) & (new_n290_ | \a[8] ) & ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))) | ((~new_n290_ ^ \a[8] ) & (~new_n291_ | ~\a[8] ) & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )))) & ((\a[5]  & ((new_n290_ & \a[8] ) | (~new_n290_ & ~\a[8] ) | ((~new_n291_ | ~\a[8] ) & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )))) & ((new_n290_ ^ \a[8] ) | (new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))) | (~\a[5]  & ((~new_n290_ ^ \a[8] ) ^ ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] ))))) | ((~\a[5]  | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )) | (new_n292_ & (~new_n291_ ^ \a[8] ))) & (new_n349_ | (\a[5]  & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )) & (~new_n292_ | (new_n291_ ^ \a[8] ))) | (~\a[5]  & (new_n292_ ^ (new_n291_ ^ \a[8] ))))))))) | (\a[5]  & ((new_n348_ & \a[8] ) | (~new_n348_ & ~\a[8] ) | ((~new_n289_ | ~\a[8] ) & ((new_n289_ & \a[8] ) | (~new_n289_ & ~\a[8] ) | ((~new_n290_ | ~\a[8] ) & ((new_n290_ & \a[8] ) | (~new_n290_ & ~\a[8] ) | ((~new_n291_ | ~\a[8] ) & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )))))))) & ((new_n348_ ^ \a[8] ) | (new_n289_ & \a[8] ) | ((~new_n289_ | ~\a[8] ) & (new_n289_ | \a[8] ) & ((new_n290_ & \a[8] ) | ((~new_n290_ | ~\a[8] ) & (new_n290_ | \a[8] ) & ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))))))) | (~\a[5]  & ((~new_n348_ ^ \a[8] ) ^ ((new_n289_ & \a[8] ) | ((~new_n289_ | ~\a[8] ) & (new_n289_ | \a[8] ) & ((new_n290_ & \a[8] ) | ((~new_n290_ | ~\a[8] ) & (new_n290_ | \a[8] ) & ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] ))))))))));
  assign new_n348_ = ~new_n214_ ^ new_n285_;
  assign new_n349_ = (~new_n350_ | ~\a[5] ) & ((new_n350_ & \a[5] ) | (~new_n350_ & ~\a[5] ) | ((~\a[5]  | ((~new_n294_ | ~\a[8] ) & (new_n294_ | \a[8] ) & ((new_n295_ & \a[8] ) | ((~new_n295_ | ~\a[8] ) & (new_n295_ | \a[8] ) & ((new_n296_ & \a[8] ) | (~new_n298_ & (~new_n296_ | ~\a[8] ) & (new_n296_ | \a[8] )))))) | ((~new_n294_ ^ \a[8] ) & (~new_n295_ | ~\a[8] ) & ((new_n295_ & \a[8] ) | (~new_n295_ & ~\a[8] ) | ((~new_n296_ | ~\a[8] ) & (new_n298_ | (new_n296_ & \a[8] ) | (~new_n296_ & ~\a[8] )))))) & ((\a[5]  & ((new_n294_ & \a[8] ) | (~new_n294_ & ~\a[8] ) | ((~new_n295_ | ~\a[8] ) & ((new_n295_ & \a[8] ) | (~new_n295_ & ~\a[8] ) | ((~new_n296_ | ~\a[8] ) & (new_n298_ | (new_n296_ & \a[8] ) | (~new_n296_ & ~\a[8] )))))) & ((new_n294_ ^ \a[8] ) | (new_n295_ & \a[8] ) | ((~new_n295_ | ~\a[8] ) & (new_n295_ | \a[8] ) & ((new_n296_ & \a[8] ) | (~new_n298_ & (~new_n296_ | ~\a[8] ) & (new_n296_ | \a[8] )))))) | (~\a[5]  & ((~new_n294_ ^ \a[8] ) ^ ((new_n295_ & \a[8] ) | ((~new_n295_ | ~\a[8] ) & (new_n295_ | \a[8] ) & ((new_n296_ & \a[8] ) | (~new_n298_ & (~new_n296_ | ~\a[8] ) & (new_n296_ | \a[8] ))))))) | ((~\a[5]  | ((~new_n295_ | ~\a[8] ) & (new_n295_ | \a[8] ) & ((new_n296_ & \a[8] ) | (~new_n298_ & (~new_n296_ | ~\a[8] ) & (new_n296_ | \a[8] )))) | ((~new_n295_ ^ \a[8] ) & (~new_n296_ | ~\a[8] ) & (new_n298_ | (new_n296_ & \a[8] ) | (~new_n296_ & ~\a[8] )))) & (new_n351_ | (\a[5]  & ((new_n295_ & \a[8] ) | (~new_n295_ & ~\a[8] ) | ((~new_n296_ | ~\a[8] ) & (new_n298_ | (new_n296_ & \a[8] ) | (~new_n296_ & ~\a[8] )))) & ((new_n295_ ^ \a[8] ) | (new_n296_ & \a[8] ) | (~new_n298_ & (~new_n296_ | ~\a[8] ) & (new_n296_ | \a[8] )))) | (~\a[5]  & ((~new_n295_ ^ \a[8] ) ^ ((new_n296_ & \a[8] ) | (~new_n298_ & (~new_n296_ | ~\a[8] ) & (new_n296_ | \a[8] ))))))))));
  assign new_n350_ = (\a[8]  ^ (~new_n219_ ^ new_n293_)) ^ ((new_n294_ & \a[8] ) | ((~new_n294_ | ~\a[8] ) & (new_n294_ | \a[8] ) & ((new_n295_ & \a[8] ) | ((~new_n295_ | ~\a[8] ) & (new_n295_ | \a[8] ) & ((new_n296_ & \a[8] ) | (~new_n298_ & (new_n296_ | \a[8] ) & (~new_n296_ | ~\a[8] )))))));
  assign new_n351_ = (~\a[5]  | (~new_n298_ & new_n352_) | (new_n298_ & ~new_n352_)) & ((\a[5]  & (new_n298_ | ~new_n352_) & (~new_n298_ | new_n352_)) | (~\a[5]  & (new_n298_ ^ new_n352_)) | ((~new_n353_ | ~\a[5] ) & ((new_n353_ & \a[5] ) | (~new_n353_ & ~\a[5] ) | ((~new_n354_ | ~\a[5] ) & ((new_n354_ & \a[5] ) | (~new_n354_ & ~\a[5] ) | ((~new_n355_ | ~\a[5] ) & (new_n356_ | (~new_n355_ & ~\a[5] ) | (new_n355_ & \a[5] ))))))));
  assign new_n352_ = \a[8]  ^ (~new_n221_ ^ new_n297_);
  assign new_n353_ = ((\a[8]  & (~new_n253_ | (~new_n226_ & (new_n229_ | ~new_n252_))) & (new_n253_ | new_n226_ | (~new_n229_ & new_n252_))) | (((~new_n334_ & (new_n229_ | ~new_n252_) & (~new_n229_ | new_n252_)) | (~new_n300_ & (new_n334_ | (~new_n229_ & new_n252_) | (new_n229_ & ~new_n252_)) & (~new_n334_ | (~new_n229_ ^ new_n252_)))) & (~\a[8]  | (new_n253_ & (new_n226_ | (~new_n229_ & new_n252_))) | (~new_n253_ & ~new_n226_ & (new_n229_ | ~new_n252_))) & (\a[8]  | (new_n253_ ^ (new_n226_ | (~new_n229_ & new_n252_)))))) ^ (new_n299_ ^ \a[8] );
  assign new_n354_ = ((~new_n334_ & (new_n229_ | ~new_n252_) & (~new_n229_ | new_n252_)) | (~new_n300_ & (new_n334_ | (~new_n229_ & new_n252_) | (new_n229_ & ~new_n252_)) & (~new_n334_ | (~new_n229_ ^ new_n252_)))) ^ (\a[8]  ^ (new_n253_ ^ (new_n226_ | (~new_n229_ & new_n252_))));
  assign new_n355_ = ~new_n300_ ^ (~new_n334_ ^ (~new_n229_ ^ new_n252_));
  assign new_n356_ = (~new_n357_ | ~\a[5] ) & (((~\a[5]  | (new_n332_ & (new_n305_ | (~new_n308_ & new_n331_))) | (~new_n332_ & ~new_n305_ & (new_n308_ | ~new_n331_))) & (((new_n391_ | (~new_n308_ & new_n331_) | (new_n308_ & ~new_n331_)) & (new_n358_ | (~new_n391_ & (new_n308_ | ~new_n331_) & (~new_n308_ | new_n331_)) | (new_n391_ & (new_n308_ ^ new_n331_)))) | (\a[5]  & (~new_n332_ | (~new_n305_ & (new_n308_ | ~new_n331_))) & (new_n332_ | new_n305_ | (~new_n308_ & new_n331_))) | (~\a[5]  & (~new_n332_ ^ (new_n305_ | (~new_n308_ & new_n331_)))))) | (new_n357_ & \a[5] ) | (~new_n357_ & ~\a[5] ));
  assign new_n357_ = (new_n303_ | (new_n332_ & (new_n305_ | (~new_n308_ & new_n331_)))) ^ (new_n301_ ^ ~new_n333_);
  assign new_n358_ = (~new_n359_ | new_n389_) & ((new_n359_ & ~new_n389_) | (~new_n359_ & new_n389_) | (~new_n361_ & (~new_n387_ | (((~new_n313_ & new_n388_) | (new_n313_ & ~new_n388_) | new_n390_) & (new_n363_ | ((new_n313_ | ~new_n388_) & (~new_n313_ | new_n388_) & ~new_n390_) | ((new_n313_ ^ new_n388_) & new_n390_))))));
  assign new_n359_ = new_n360_ ^ (new_n311_ | (new_n327_ & ((~new_n330_ & (new_n240_ | (~new_n239_ & new_n247_) | (new_n239_ & ~new_n247_)) & (~new_n240_ | (~new_n239_ ^ new_n247_))) | (~new_n313_ & (new_n330_ | (~new_n240_ & (new_n239_ | ~new_n247_) & (~new_n239_ | new_n247_)) | (new_n240_ & (new_n239_ ^ new_n247_))) & (~new_n330_ | (~new_n240_ ^ (~new_n239_ ^ new_n247_)))))));
  assign new_n360_ = ~new_n328_ ^ ((~new_n235_ ^ new_n236_) ^ ((new_n237_ & ~new_n238_) | ((new_n237_ | ~new_n238_) & (~new_n237_ | new_n238_) & ((~new_n239_ & new_n247_) | (~new_n240_ & (new_n239_ | ~new_n247_) & (~new_n239_ | new_n247_))))));
  assign new_n361_ = ~new_n362_ & (~new_n327_ | ((new_n330_ | (~new_n240_ & (new_n239_ | ~new_n247_) & (~new_n239_ | new_n247_)) | (new_n240_ & (new_n239_ ^ new_n247_))) & (new_n313_ | (~new_n330_ & (new_n240_ | (~new_n239_ & new_n247_) | (new_n239_ & ~new_n247_)) & (~new_n240_ | (~new_n239_ ^ new_n247_))) | (new_n330_ & (new_n240_ ^ (~new_n239_ ^ new_n247_)))))) & (new_n327_ | (~new_n330_ & (new_n240_ | (~new_n239_ & new_n247_) | (new_n239_ & ~new_n247_)) & (~new_n240_ | (~new_n239_ ^ new_n247_))) | (~new_n313_ & (new_n330_ | (~new_n240_ & (new_n239_ | ~new_n247_) & (~new_n239_ | new_n247_)) | (new_n240_ & (new_n239_ ^ new_n247_))) & (~new_n330_ | (~new_n240_ ^ (~new_n239_ ^ new_n247_)))));
  assign new_n362_ = \a[5]  ^ ((~new_n116_ | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[11]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[12]  | (~\a[4]  ^ ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[10]  | (~\a[3]  ^ ~\a[4] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n363_ = (~new_n365_ | new_n384_) & ((new_n365_ & ~new_n384_) | (~new_n365_ & new_n384_) | (~new_n366_ & (~new_n368_ | ((new_n386_ | (new_n364_ & ~new_n319_) | (~new_n364_ & new_n319_)) & (new_n369_ | (~new_n386_ & (~new_n364_ | new_n319_) & (new_n364_ | ~new_n319_)) | (new_n386_ & (~new_n364_ ^ ~new_n319_)))))));
  assign new_n364_ = ~new_n318_ ^ new_n326_;
  assign new_n365_ = (~new_n314_ ^ new_n315_) ^ ((new_n316_ & ~new_n317_) | (((~new_n318_ & new_n326_) | (~new_n319_ & (new_n318_ | ~new_n326_) & (~new_n318_ | new_n326_))) & (new_n316_ | ~new_n317_) & (~new_n316_ | new_n317_)));
  assign new_n366_ = ~new_n367_ & ((~new_n316_ & new_n317_) | (new_n316_ & ~new_n317_) | ((new_n318_ | ~new_n326_) & (new_n319_ | (~new_n318_ & new_n326_) | (new_n318_ & ~new_n326_)))) & ((~new_n316_ ^ new_n317_) | (~new_n318_ & new_n326_) | (~new_n319_ & (new_n318_ | ~new_n326_) & (~new_n318_ | new_n326_)));
  assign new_n367_ = \a[5]  ^ (((~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n73_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[9]  | (~\a[4]  ^ ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[7]  | (~\a[3]  ^ ~\a[4] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n368_ = ~new_n367_ ^ ((~new_n316_ ^ new_n317_) ^ ((~new_n318_ & new_n326_) | (~new_n319_ & (new_n318_ | ~new_n326_) & (~new_n318_ | new_n326_))));
  assign new_n369_ = (~new_n370_ | new_n371_) & ((~new_n370_ & new_n371_) | (new_n370_ & ~new_n371_) | ((~new_n372_ | new_n373_) & (((new_n374_ | ~new_n383_) & (new_n377_ | (~new_n374_ & new_n383_) | (new_n374_ & ~new_n383_))) | (~new_n372_ & new_n373_) | (new_n372_ & ~new_n373_))));
  assign new_n370_ = (new_n323_ | (~new_n324_ & new_n325_)) ^ (new_n322_ ^ (~\a[8]  ^ (new_n321_ & (~new_n63_ | ~new_n320_))));
  assign new_n371_ = \a[5]  ^ ((~new_n54_ | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[6]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[7]  | (~\a[4]  ^ ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[5]  | (~\a[3]  ^ ~\a[4] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n372_ = ~new_n324_ ^ new_n325_;
  assign new_n373_ = \a[5]  ^ ((~new_n57_ | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[5]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[6]  | (~\a[4]  ^ ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[4]  | (~\a[3]  ^ ~\a[4] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n374_ = \a[5]  ^ (new_n376_ & (~new_n60_ | ~new_n375_));
  assign new_n375_ = (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (\a[4]  | \a[5] ) & (~\a[4]  | ~\a[5] );
  assign new_n376_ = (~\b[4]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[5]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[3]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n377_ = (~new_n379_ | (\a[5]  ^ (new_n378_ & (~new_n63_ | ~new_n375_)))) & ((~new_n380_ & (new_n381_ | ~new_n382_)) | (new_n379_ & (~\a[5]  ^ (new_n378_ & (~new_n63_ | ~new_n375_)))) | (~new_n379_ & (~\a[5]  | ~new_n378_ | (new_n63_ & new_n375_)) & (\a[5]  | (new_n378_ & (~new_n63_ | ~new_n375_)))));
  assign new_n378_ = (~\b[3]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[4]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[2]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n379_ = ((\b[0]  & (\a[5]  ^ ~\a[6] ) & (\a[6]  | \a[7] ) & (~\a[6]  | ~\a[7] )) | (\b[1]  & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (\a[7]  ^ ~\a[8] )) | ((\b[0]  ^ \b[1] ) & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] ))) ^ (\a[8]  & \b[0]  & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ));
  assign new_n380_ = \b[0]  & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (~\b[0]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\b[0]  ^ \b[1] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[1]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n381_ = \a[5]  ^ (((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[2]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )));
  assign new_n382_ = (\b[0]  & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] )) ^ ((~\b[0]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\b[0]  ^ \b[1] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[1]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )));
  assign new_n383_ = (~\a[8]  | ((~\b[0]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\b[0]  ^ \b[1] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )))) ^ ((~\b[1]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[2]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )));
  assign new_n384_ = \a[5]  ^ (new_n385_ & (~new_n375_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n73_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n385_ = (~\b[9]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[10]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[8]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n386_ = \a[5]  ^ (((~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n73_ & (~\b[7]  ^ \b[8] ))) & (~\b[7]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[8]  | (~\a[4]  ^ ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[6]  | (~\a[3]  ^ ~\a[4] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n387_ = ~new_n362_ ^ (new_n327_ ^ ((~new_n330_ & (new_n240_ | (~new_n239_ & new_n247_) | (new_n239_ & ~new_n247_)) & (~new_n240_ | (~new_n239_ ^ new_n247_))) | (~new_n313_ & (new_n330_ | (~new_n240_ & (new_n239_ | ~new_n247_) & (~new_n239_ | new_n247_)) | (new_n240_ & (new_n239_ ^ new_n247_))) & (~new_n330_ | (~new_n240_ ^ (~new_n239_ ^ new_n247_))))));
  assign new_n388_ = ~new_n330_ ^ (~new_n240_ ^ (~new_n239_ ^ new_n247_));
  assign new_n389_ = \a[5]  ^ (((new_n82_ ^ \b[12] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[12]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[11]  | (~\a[3]  ^ ~\a[4] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n390_ = \a[5]  ^ ((~new_n89_ | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[10]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[11]  | (~\a[4]  ^ ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[9]  | (~\a[3]  ^ ~\a[4] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n391_ = \a[5]  ^ (~\b[12]  | ((new_n82_ | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[3]  ^ ~\a[4] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  ^ ~\a[3] ))));
  assign new_n392_ = \a[5]  ^ (~new_n286_ ^ (new_n283_ ^ \a[8] ));
  assign new_n393_ = (new_n342_ ^ \a[5] ) ^ ((new_n343_ & \a[5] ) | ((new_n344_ | (~new_n345_ & new_n392_)) & (~new_n343_ | ~\a[5] ) & (new_n343_ | \a[5] )));
  assign new_n394_ = (new_n343_ ^ \a[5] ) ^ (new_n344_ | (~new_n345_ & new_n392_));
  assign new_n395_ = (~\a[2]  | (new_n396_ & ~new_n347_) | (~new_n396_ & new_n347_)) & (((~new_n445_ | ~\a[2] ) & ((~new_n445_ & ~\a[2] ) | (new_n445_ & \a[2] ) | ((~new_n446_ | ~\a[2] ) & (new_n397_ | (new_n446_ & \a[2] ) | (~new_n446_ & ~\a[2] ))))) | (\a[2]  & (~new_n396_ | new_n347_) & (new_n396_ | ~new_n347_)) | (~\a[2]  & (~new_n396_ ^ ~new_n347_)));
  assign new_n396_ = ~new_n346_ ^ ~\a[5] ;
  assign new_n397_ = (~\a[2]  | (((\a[5]  & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )) & (~new_n292_ | (new_n291_ ^ \a[8] ))) | (~new_n349_ & (~\a[5]  | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )) | (new_n292_ & (~new_n291_ ^ \a[8] ))) & (\a[5]  | (~new_n292_ ^ (new_n291_ ^ \a[8] ))))) & (~\a[5]  | ((~new_n290_ | ~\a[8] ) & (new_n290_ | \a[8] ) & ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))) | ((~new_n290_ ^ \a[8] ) & (~new_n291_ | ~\a[8] ) & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )))) & (\a[5]  | ((new_n290_ ^ \a[8] ) ^ ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))))) | ((~\a[5]  | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )) | (new_n292_ & (~new_n291_ ^ \a[8] ))) & (new_n349_ | (\a[5]  & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )) & (~new_n292_ | (new_n291_ ^ \a[8] ))) | (~\a[5]  & (new_n292_ ^ (new_n291_ ^ \a[8] )))) & (~\a[5]  ^ ((new_n290_ ^ \a[8] ) ^ ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] ))))))) & (new_n398_ | (\a[2]  & (((~\a[5]  | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )) | (new_n292_ & (~new_n291_ ^ \a[8] ))) & (new_n349_ | (\a[5]  & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )) & (~new_n292_ | (new_n291_ ^ \a[8] ))) | (~\a[5]  & (new_n292_ ^ (new_n291_ ^ \a[8] ))))) | (\a[5]  & ((new_n290_ & \a[8] ) | (~new_n290_ & ~\a[8] ) | ((~new_n291_ | ~\a[8] ) & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )))) & ((new_n290_ ^ \a[8] ) | (new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))) | (~\a[5]  & ((~new_n290_ ^ \a[8] ) ^ ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))))) & ((\a[5]  & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )) & (~new_n292_ | (new_n291_ ^ \a[8] ))) | (~new_n349_ & (~\a[5]  | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )) | (new_n292_ & (~new_n291_ ^ \a[8] ))) & (\a[5]  | (~new_n292_ ^ (new_n291_ ^ \a[8] )))) | (\a[5]  ^ ((new_n290_ ^ \a[8] ) ^ ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] ))))))) | (~\a[2]  & (((~\a[5]  | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )) | (new_n292_ & (~new_n291_ ^ \a[8] ))) & (new_n349_ | (\a[5]  & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )) & (~new_n292_ | (new_n291_ ^ \a[8] ))) | (~\a[5]  & (new_n292_ ^ (new_n291_ ^ \a[8] ))))) ^ (\a[5]  ^ ((new_n290_ ^ \a[8] ) ^ ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] ))))))));
  assign new_n398_ = (~\a[2]  | (new_n401_ & ((new_n350_ & \a[5] ) | (~new_n399_ & (new_n350_ | \a[5] ) & (~new_n350_ | ~\a[5] )))) | (~new_n401_ & (~new_n350_ | ~\a[5] ) & (new_n399_ | (~new_n350_ & ~\a[5] ) | (new_n350_ & \a[5] )))) & (((~\a[2]  | (~new_n399_ & (new_n350_ | \a[5] ) & (~new_n350_ | ~\a[5] )) | (new_n399_ & (new_n350_ ^ ~\a[5] ))) & (((~new_n402_ | ~\a[2] ) & (new_n403_ | (~new_n402_ & ~\a[2] ) | (new_n402_ & \a[2] ))) | (\a[2]  & (new_n399_ | (~new_n350_ & ~\a[5] ) | (new_n350_ & \a[5] )) & (~new_n399_ | (~new_n350_ ^ ~\a[5] ))) | (~\a[2]  & (new_n399_ ^ (~new_n350_ ^ ~\a[5] ))))) | (\a[2]  & (~new_n401_ | ((~new_n350_ | ~\a[5] ) & (new_n399_ | (~new_n350_ & ~\a[5] ) | (new_n350_ & \a[5] )))) & (new_n401_ | (new_n350_ & \a[5] ) | (~new_n399_ & (new_n350_ | \a[5] ) & (~new_n350_ | ~\a[5] )))) | (~\a[2]  & (~new_n401_ ^ ((new_n350_ & \a[5] ) | (~new_n399_ & (new_n350_ | \a[5] ) & (~new_n350_ | ~\a[5] ))))));
  assign new_n399_ = (~\a[5]  | ((~new_n294_ | ~\a[8] ) & (new_n294_ | \a[8] ) & ((new_n295_ & \a[8] ) | ((~new_n295_ | ~\a[8] ) & (new_n295_ | \a[8] ) & ((~new_n298_ & new_n352_) | (new_n296_ & \a[8] ))))) | ((~new_n294_ ^ \a[8] ) & (~new_n295_ | ~\a[8] ) & ((new_n295_ & \a[8] ) | (~new_n295_ & ~\a[8] ) | ((new_n298_ | ~new_n352_) & (~new_n296_ | ~\a[8] ))))) & (((~\a[5]  | ((~new_n295_ | ~\a[8] ) & (new_n295_ | \a[8] ) & ((~new_n298_ & new_n352_) | (new_n296_ & \a[8] ))) | ((~new_n295_ ^ \a[8] ) & (new_n298_ | ~new_n352_) & (~new_n296_ | ~\a[8] ))) & (((~\a[5]  | (~new_n298_ & new_n352_) | (new_n298_ & ~new_n352_)) & (new_n400_ | (\a[5]  & (new_n298_ | ~new_n352_) & (~new_n298_ | new_n352_)) | (~\a[5]  & (new_n298_ ^ new_n352_)))) | (\a[5]  & ((new_n295_ & \a[8] ) | (~new_n295_ & ~\a[8] ) | ((new_n298_ | ~new_n352_) & (~new_n296_ | ~\a[8] ))) & ((new_n295_ ^ \a[8] ) | (~new_n298_ & new_n352_) | (new_n296_ & \a[8] ))) | (~\a[5]  & ((~new_n295_ ^ \a[8] ) ^ ((~new_n298_ & new_n352_) | (new_n296_ & \a[8] )))))) | (\a[5]  & ((new_n294_ & \a[8] ) | (~new_n294_ & ~\a[8] ) | ((~new_n295_ | ~\a[8] ) & ((new_n295_ & \a[8] ) | (~new_n295_ & ~\a[8] ) | ((new_n298_ | ~new_n352_) & (~new_n296_ | ~\a[8] ))))) & ((new_n294_ ^ \a[8] ) | (new_n295_ & \a[8] ) | ((~new_n295_ | ~\a[8] ) & (new_n295_ | \a[8] ) & ((~new_n298_ & new_n352_) | (new_n296_ & \a[8] ))))) | (~\a[5]  & ((~new_n294_ ^ \a[8] ) ^ ((new_n295_ & \a[8] ) | ((~new_n295_ | ~\a[8] ) & (new_n295_ | \a[8] ) & ((~new_n298_ & new_n352_) | (new_n296_ & \a[8] )))))));
  assign new_n400_ = (~new_n353_ | ~\a[5] ) & ((new_n353_ & \a[5] ) | (~new_n353_ & ~\a[5] ) | ((~new_n354_ | ~\a[5] ) & ((~new_n354_ & ~\a[5] ) | (new_n354_ & \a[5] ) | ((~new_n355_ | ~\a[5] ) & (new_n356_ | (new_n355_ & \a[5] ) | (~new_n355_ & ~\a[5] ))))));
  assign new_n401_ = \a[5]  ^ (~new_n292_ ^ (new_n291_ ^ \a[8] ));
  assign new_n402_ = ((\a[5]  & ((new_n295_ & \a[8] ) | (~new_n295_ & ~\a[8] ) | ((new_n298_ | ~new_n352_) & (~new_n296_ | ~\a[8] ))) & ((new_n295_ ^ \a[8] ) | (~new_n298_ & new_n352_) | (new_n296_ & \a[8] ))) | (((\a[5]  & (new_n298_ | ~new_n352_) & (~new_n298_ | new_n352_)) | (~new_n400_ & (~\a[5]  | (~new_n298_ & new_n352_) | (new_n298_ & ~new_n352_)) & (\a[5]  | (~new_n298_ ^ new_n352_)))) & (~\a[5]  | ((~new_n295_ | ~\a[8] ) & (new_n295_ | \a[8] ) & ((~new_n298_ & new_n352_) | (new_n296_ & \a[8] ))) | ((~new_n295_ ^ \a[8] ) & (new_n298_ | ~new_n352_) & (~new_n296_ | ~\a[8] ))) & (\a[5]  | ((new_n295_ ^ \a[8] ) ^ ((~new_n298_ & new_n352_) | (new_n296_ & \a[8] )))))) ^ (\a[5]  ^ ((new_n294_ ^ \a[8] ) ^ ((new_n295_ & \a[8] ) | ((~new_n295_ | ~\a[8] ) & (new_n295_ | \a[8] ) & ((~new_n298_ & new_n352_) | (new_n296_ & \a[8] ))))));
  assign new_n403_ = (~\a[2]  | (new_n404_ & (((new_n298_ | ~new_n352_) & (~new_n298_ | new_n352_) & \a[5] ) | (~new_n400_ & ((~new_n298_ & new_n352_) | (new_n298_ & ~new_n352_) | ~\a[5] ) & ((~new_n298_ ^ new_n352_) | \a[5] )))) | (~new_n404_ & ((~new_n298_ & new_n352_) | (new_n298_ & ~new_n352_) | ~\a[5] ) & (new_n400_ | ((new_n298_ | ~new_n352_) & (~new_n298_ | new_n352_) & \a[5] ) | ((new_n298_ ^ new_n352_) & ~\a[5] )))) & (((~\a[2]  | (~new_n400_ & ((~new_n298_ & new_n352_) | (new_n298_ & ~new_n352_) | ~\a[5] ) & ((~new_n298_ ^ new_n352_) | \a[5] )) | (new_n400_ & ((new_n298_ ^ new_n352_) ^ \a[5] ))) & (((~new_n405_ | ~\a[2] ) & (new_n406_ | (new_n405_ & \a[2] ) | (~new_n405_ & ~\a[2] ))) | (\a[2]  & (new_n400_ | ((new_n298_ | ~new_n352_) & (~new_n298_ | new_n352_) & \a[5] ) | ((new_n298_ ^ new_n352_) & ~\a[5] )) & (~new_n400_ | ((~new_n298_ ^ new_n352_) ^ \a[5] ))) | (~\a[2]  & (new_n400_ ^ ((~new_n298_ ^ new_n352_) ^ \a[5] ))))) | (\a[2]  & (~new_n404_ | (((~new_n298_ & new_n352_) | (new_n298_ & ~new_n352_) | ~\a[5] ) & (new_n400_ | ((new_n298_ | ~new_n352_) & (~new_n298_ | new_n352_) & \a[5] ) | ((new_n298_ ^ new_n352_) & ~\a[5] )))) & (new_n404_ | ((new_n298_ | ~new_n352_) & (~new_n298_ | new_n352_) & \a[5] ) | (~new_n400_ & ((~new_n298_ & new_n352_) | (new_n298_ & ~new_n352_) | ~\a[5] ) & ((~new_n298_ ^ new_n352_) | \a[5] )))) | (~\a[2]  & (~new_n404_ ^ (((new_n298_ | ~new_n352_) & (~new_n298_ | new_n352_) & \a[5] ) | (~new_n400_ & ((~new_n298_ & new_n352_) | (new_n298_ & ~new_n352_) | ~\a[5] ) & ((~new_n298_ ^ new_n352_) | \a[5] ))))));
  assign new_n404_ = \a[5]  ^ ((new_n295_ ^ \a[8] ) ^ ((new_n296_ & \a[8] ) | (~new_n298_ & (new_n296_ | \a[8] ) & (~new_n296_ | ~\a[8] ))));
  assign new_n405_ = (new_n353_ ^ \a[5] ) ^ ((new_n354_ & \a[5] ) | ((new_n354_ | \a[5] ) & (~new_n354_ | ~\a[5] ) & ((new_n355_ & \a[5] ) | (~new_n356_ & (~new_n355_ | ~\a[5] ) & (new_n355_ | \a[5] )))));
  assign new_n406_ = (~\a[2]  | ((~new_n354_ | ~\a[5] ) & (new_n354_ | \a[5] ) & ((new_n355_ & \a[5] ) | (~new_n356_ & (~new_n355_ | ~\a[5] ) & (new_n355_ | \a[5] )))) | ((~new_n354_ ^ \a[5] ) & (~new_n355_ | ~\a[5] ) & (new_n356_ | (new_n355_ & \a[5] ) | (~new_n355_ & ~\a[5] )))) & (((~\a[2]  | (~new_n356_ & (~new_n355_ | ~\a[5] ) & (new_n355_ | \a[5] )) | (new_n356_ & (~new_n355_ ^ \a[5] ))) & (((~new_n407_ | ~\a[2] ) & ((new_n407_ & \a[2] ) | (~new_n407_ & ~\a[2] ) | ((~new_n408_ | ~\a[2] ) & (new_n409_ | (~new_n408_ & ~\a[2] ) | (new_n408_ & \a[2] ))))) | (\a[2]  & (new_n356_ | (new_n355_ & \a[5] ) | (~new_n355_ & ~\a[5] )) & (~new_n356_ | (new_n355_ ^ \a[5] ))) | (~\a[2]  & (new_n356_ ^ (new_n355_ ^ \a[5] ))))) | (\a[2]  & ((new_n354_ & \a[5] ) | (~new_n354_ & ~\a[5] ) | ((~new_n355_ | ~\a[5] ) & (new_n356_ | (new_n355_ & \a[5] ) | (~new_n355_ & ~\a[5] )))) & ((new_n354_ ^ \a[5] ) | (new_n355_ & \a[5] ) | (~new_n356_ & (~new_n355_ | ~\a[5] ) & (new_n355_ | \a[5] )))) | (~\a[2]  & ((~new_n354_ ^ \a[5] ) ^ ((new_n355_ & \a[5] ) | (~new_n356_ & (~new_n355_ | ~\a[5] ) & (new_n355_ | \a[5] ))))));
  assign new_n407_ = ((\a[5]  & (~new_n332_ | (~new_n305_ & (new_n308_ | ~new_n331_))) & (new_n332_ | new_n305_ | (~new_n308_ & new_n331_))) | (((~new_n391_ & (new_n308_ | ~new_n331_) & (~new_n308_ | new_n331_)) | (~new_n358_ & (new_n391_ | (~new_n308_ & new_n331_) | (new_n308_ & ~new_n331_)) & (~new_n391_ | (~new_n308_ ^ new_n331_)))) & (~\a[5]  | (new_n332_ & (new_n305_ | (~new_n308_ & new_n331_))) | (~new_n332_ & ~new_n305_ & (new_n308_ | ~new_n331_))) & (\a[5]  | (new_n332_ ^ (new_n305_ | (~new_n308_ & new_n331_)))))) ^ (new_n357_ ^ \a[5] );
  assign new_n408_ = ((~new_n391_ & (new_n308_ | ~new_n331_) & (~new_n308_ | new_n331_)) | (~new_n358_ & (new_n391_ | (~new_n308_ & new_n331_) | (new_n308_ & ~new_n331_)) & (~new_n391_ | (~new_n308_ ^ new_n331_)))) ^ (\a[5]  ^ (new_n332_ ^ (new_n305_ | (~new_n308_ & new_n331_))));
  assign new_n409_ = (~\a[2]  | (~new_n358_ & new_n410_) | (new_n358_ & ~new_n410_)) & ((\a[2]  & (new_n358_ | ~new_n410_) & (~new_n358_ | new_n410_)) | (~\a[2]  & (new_n358_ ^ new_n410_)) | ((~new_n411_ | ~\a[2] ) & ((new_n411_ & \a[2] ) | (~new_n411_ & ~\a[2] ) | (~new_n412_ & (new_n413_ | ~new_n444_)))));
  assign new_n410_ = ~new_n391_ ^ (~new_n308_ ^ new_n331_);
  assign new_n411_ = (new_n359_ ^ ~new_n389_) ^ (new_n361_ | (new_n387_ & (((new_n313_ | ~new_n388_) & (~new_n313_ | new_n388_) & ~new_n390_) | (~new_n363_ & ((~new_n313_ & new_n388_) | (new_n313_ & ~new_n388_) | new_n390_) & ((~new_n313_ ^ new_n388_) | ~new_n390_)))));
  assign new_n412_ = \a[2]  & (~new_n387_ | ((new_n390_ | (~new_n313_ & new_n388_) | (new_n313_ & ~new_n388_)) & (new_n363_ | (~new_n390_ & (new_n313_ | ~new_n388_) & (~new_n313_ | new_n388_)) | (new_n390_ & (new_n313_ ^ new_n388_))))) & (new_n387_ | (~new_n390_ & (new_n313_ | ~new_n388_) & (~new_n313_ | new_n388_)) | (~new_n363_ & (new_n390_ | (~new_n313_ & new_n388_) | (new_n313_ & ~new_n388_)) & (~new_n390_ | (~new_n313_ ^ new_n388_))));
  assign new_n413_ = (new_n442_ | (~new_n363_ & new_n414_) | (new_n363_ & ~new_n414_)) & (((~new_n415_ | new_n443_) & ((~new_n417_ & (new_n419_ | ~new_n441_)) | (new_n415_ & ~new_n443_) | (~new_n415_ & new_n443_))) | (~new_n442_ & (new_n363_ | ~new_n414_) & (~new_n363_ | new_n414_)) | (new_n442_ & (new_n363_ ^ new_n414_)));
  assign new_n414_ = ~new_n390_ ^ (~new_n313_ ^ new_n388_);
  assign new_n415_ = new_n416_ ^ (new_n366_ | (new_n368_ & ((~new_n386_ & (new_n319_ | (~new_n318_ & new_n326_) | (new_n318_ & ~new_n326_)) & (~new_n319_ | (~new_n318_ ^ new_n326_))) | (~new_n369_ & (new_n386_ | (~new_n319_ & (new_n318_ | ~new_n326_) & (~new_n318_ | new_n326_)) | (new_n319_ & (new_n318_ ^ new_n326_))) & (~new_n386_ | (~new_n319_ ^ (~new_n318_ ^ new_n326_)))))));
  assign new_n416_ = ~new_n384_ ^ ((~new_n314_ ^ new_n315_) ^ ((new_n316_ & ~new_n317_) | ((new_n316_ | ~new_n317_) & (~new_n316_ | new_n317_) & ((~new_n318_ & new_n326_) | (~new_n319_ & (new_n318_ | ~new_n326_) & (~new_n318_ | new_n326_))))));
  assign new_n417_ = ~new_n418_ & (~new_n368_ | ((new_n386_ | (~new_n319_ & (new_n318_ | ~new_n326_) & (~new_n318_ | new_n326_)) | (new_n319_ & (new_n318_ ^ new_n326_))) & (new_n369_ | (~new_n386_ & (new_n319_ | (~new_n318_ & new_n326_) | (new_n318_ & ~new_n326_)) & (~new_n319_ | (~new_n318_ ^ new_n326_))) | (new_n386_ & (new_n319_ ^ (~new_n318_ ^ new_n326_)))))) & (new_n368_ | (~new_n386_ & (new_n319_ | (~new_n318_ & new_n326_) | (new_n318_ & ~new_n326_)) & (~new_n319_ | (~new_n318_ ^ new_n326_))) | (~new_n369_ & (new_n386_ | (~new_n319_ & (new_n318_ | ~new_n326_) & (~new_n318_ | new_n326_)) | (new_n319_ & (new_n318_ ^ new_n326_))) & (~new_n386_ | (~new_n319_ ^ (~new_n318_ ^ new_n326_)))));
  assign new_n418_ = \a[2]  ^ ((~new_n116_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[10]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[12]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[11]  | \a[0]  | ~\a[1] ));
  assign new_n419_ = (new_n421_ | (~new_n369_ & new_n420_) | (new_n369_ & ~new_n420_)) & ((~new_n421_ & (new_n369_ | ~new_n420_) & (~new_n369_ | new_n420_)) | (new_n421_ & (new_n369_ ^ new_n420_)) | ((~new_n422_ | new_n440_) & ((~new_n423_ & (new_n425_ | ~new_n439_)) | (new_n422_ & ~new_n440_) | (~new_n422_ & new_n440_))));
  assign new_n420_ = ~new_n386_ ^ (~new_n319_ ^ (~new_n318_ ^ new_n326_));
  assign new_n421_ = \a[2]  ^ ((~new_n89_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[9]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[11]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[10]  | \a[0]  | ~\a[1] ));
  assign new_n422_ = (~new_n370_ ^ new_n371_) ^ ((new_n372_ & ~new_n373_) | (((~new_n374_ & new_n383_) | (~new_n377_ & (new_n374_ | ~new_n383_) & (~new_n374_ | new_n383_))) & (new_n372_ | ~new_n373_) & (~new_n372_ | new_n373_)));
  assign new_n423_ = ~new_n424_ & ((~new_n372_ & new_n373_) | (new_n372_ & ~new_n373_) | ((new_n374_ | ~new_n383_) & (new_n377_ | (~new_n374_ & new_n383_) | (new_n374_ & ~new_n383_)))) & ((~new_n372_ ^ new_n373_) | (~new_n374_ & new_n383_) | (~new_n377_ & (new_n374_ | ~new_n383_) & (~new_n374_ | new_n383_)));
  assign new_n424_ = \a[2]  ^ ((~\b[7]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[9]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[8]  | \a[0]  | ~\a[1] ) & (~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n73_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))));
  assign new_n425_ = (new_n427_ | (~new_n377_ & new_n426_) | (new_n377_ & ~new_n426_)) & ((~new_n427_ & (new_n377_ | ~new_n426_) & (~new_n377_ | new_n426_)) | (new_n427_ & (new_n377_ ^ new_n426_)) | ((new_n428_ | ~new_n429_) & ((~new_n428_ & new_n429_) | (new_n428_ & ~new_n429_) | ((new_n430_ | ~new_n431_) & (new_n432_ | (~new_n430_ & new_n431_) | (new_n430_ & ~new_n431_))))));
  assign new_n426_ = new_n383_ ^ (~\a[5]  ^ (new_n376_ & (~new_n60_ | ~new_n375_)));
  assign new_n427_ = \a[2]  ^ ((~\b[6]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[8]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[7]  | \a[0]  | ~\a[1] ) & (~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n73_ & (~\b[7]  ^ \b[8] ))));
  assign new_n428_ = \a[2]  ^ ((~new_n54_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[5]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[7]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[6]  | \a[0]  | ~\a[1] ));
  assign new_n429_ = (new_n380_ | (~new_n381_ & new_n382_)) ^ (new_n379_ ^ (~\a[5]  ^ (new_n378_ & (~new_n63_ | ~new_n375_))));
  assign new_n430_ = \a[2]  ^ ((~new_n57_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[4]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[6]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[5]  | \a[0]  | ~\a[1] ));
  assign new_n431_ = ~new_n381_ ^ new_n382_;
  assign new_n432_ = (~new_n435_ | (\a[2]  ^ (new_n434_ & (~new_n60_ | ~new_n433_)))) & ((new_n435_ & (~\a[2]  ^ (new_n434_ & (~new_n60_ | ~new_n433_)))) | (~new_n435_ & (~\a[2]  | ~new_n434_ | (new_n60_ & new_n433_)) & (\a[2]  | (new_n434_ & (~new_n60_ | ~new_n433_)))) | ((new_n436_ | ~new_n437_) & (~new_n438_ | (~new_n436_ & new_n437_) | (new_n436_ & ~new_n437_))));
  assign new_n433_ = \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] );
  assign new_n434_ = (~\b[3]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[5]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[4]  | \a[0]  | ~\a[1] );
  assign new_n435_ = (~\a[5]  | ((~\b[0]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\b[0]  ^ \b[1] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )))) ^ ((~\b[1]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[2]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )));
  assign new_n436_ = \a[2]  ^ ((~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )))) | ((~\b[3]  ^ \b[4] ) & (~\b[2]  | ~\b[3] ) & ((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[4]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[3]  | \a[0]  | ~\a[1] ));
  assign new_n437_ = ((\b[0]  & (\a[2]  ^ ~\a[3] ) & (\a[3]  | \a[4] ) & (~\a[3]  | ~\a[4] )) | (\b[1]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (\a[4]  ^ ~\a[5] )) | ((\b[0]  ^ \b[1] ) & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (\a[4]  | \a[5] ) & (~\a[4]  | ~\a[5] ))) ^ (\a[5]  & \b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ));
  assign new_n438_ = ((\b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] )) | (\a[2]  & (~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] ) & (((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))) | (~\a[2]  & ((\b[1]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[3]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[2]  & ~\a[0]  & \a[1] ) | (((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )) & ((\b[2]  ^ \b[3] ) | (\b[1]  & (\b[0]  | \b[2] ))) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] ))))) & ((\b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (~\a[2]  ^ ((~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] ) & (((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))))) | ((~\b[2]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[1]  | \a[0]  | ~\a[1] ) & (~\b[0]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & ((\b[2]  ^ (\b[0]  | ~\b[1] )) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[0]  | \a[0]  | ~\a[1] ) & (~\b[1]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & ((~\b[0]  ^ \b[1] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & \a[2]  & (~\a[0]  | ~\b[0] )));
  assign new_n439_ = ~new_n424_ ^ ((~new_n372_ ^ new_n373_) ^ ((~new_n374_ & new_n383_) | (~new_n377_ & (new_n374_ | ~new_n383_) & (~new_n374_ | new_n383_))));
  assign new_n440_ = \a[2]  ^ ((((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n73_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n73_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[8]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[10]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[9]  | \a[0]  | ~\a[1] ));
  assign new_n441_ = ~new_n418_ ^ (new_n368_ ^ ((~new_n386_ & (new_n319_ | (~new_n318_ & new_n326_) | (new_n318_ & ~new_n326_)) & (~new_n319_ | (~new_n318_ ^ new_n326_))) | (~new_n369_ & (new_n386_ | (~new_n319_ & (new_n318_ | ~new_n326_) & (~new_n318_ | new_n326_)) | (new_n319_ & (new_n318_ ^ new_n326_))) & (~new_n386_ | (~new_n319_ ^ (~new_n318_ ^ new_n326_))))));
  assign new_n442_ = \a[2]  ^ (~\b[12]  | (((~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (new_n82_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))));
  assign new_n443_ = \a[2]  ^ (((new_n82_ ^ \b[12] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[11]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[12]  | \a[0]  | ~\a[1] ));
  assign new_n444_ = \a[2]  ^ (new_n387_ ^ ((~new_n390_ & (new_n313_ | ~new_n388_) & (~new_n313_ | new_n388_)) | (~new_n363_ & (new_n390_ | (~new_n313_ & new_n388_) | (new_n313_ & ~new_n388_)) & (~new_n390_ | (~new_n313_ ^ new_n388_)))));
  assign new_n445_ = ((\a[5]  & ((new_n289_ & \a[8] ) | (~new_n289_ & ~\a[8] ) | ((~new_n290_ | ~\a[8] ) & ((new_n290_ & \a[8] ) | (~new_n290_ & ~\a[8] ) | ((~new_n291_ | ~\a[8] ) & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )))))) & ((new_n289_ ^ \a[8] ) | (new_n290_ & \a[8] ) | ((~new_n290_ | ~\a[8] ) & (new_n290_ | \a[8] ) & ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))))) | ((~\a[5]  | ((~new_n289_ | ~\a[8] ) & (new_n289_ | \a[8] ) & ((new_n290_ & \a[8] ) | ((~new_n290_ | ~\a[8] ) & (new_n290_ | \a[8] ) & ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))))) | ((~new_n289_ ^ \a[8] ) & (~new_n290_ | ~\a[8] ) & ((new_n290_ & \a[8] ) | (~new_n290_ & ~\a[8] ) | ((~new_n291_ | ~\a[8] ) & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )))))) & (\a[5]  | ((new_n289_ ^ \a[8] ) ^ ((new_n290_ & \a[8] ) | ((~new_n290_ | ~\a[8] ) & (new_n290_ | \a[8] ) & ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] ))))))) & ((\a[5]  & ((new_n290_ & \a[8] ) | (~new_n290_ & ~\a[8] ) | ((~new_n291_ | ~\a[8] ) & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )))) & ((new_n290_ ^ \a[8] ) | (new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))) | ((~\a[5]  | ((~new_n290_ | ~\a[8] ) & (new_n290_ | \a[8] ) & ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))) | ((~new_n290_ ^ \a[8] ) & (~new_n291_ | ~\a[8] ) & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )))) & (\a[5]  | ((new_n290_ ^ \a[8] ) ^ ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] ))))) & ((\a[5]  & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )) & (~new_n292_ | (new_n291_ ^ \a[8] ))) | (~new_n349_ & (~\a[5]  | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )) | (new_n292_ & (~new_n291_ ^ \a[8] ))) & (\a[5]  | (~new_n292_ ^ (new_n291_ ^ \a[8] ))))))))) ^ (\a[5]  ^ ((new_n348_ ^ \a[8] ) ^ ((new_n289_ & \a[8] ) | ((~new_n289_ | ~\a[8] ) & (new_n289_ | \a[8] ) & ((new_n290_ & \a[8] ) | ((~new_n290_ | ~\a[8] ) & (new_n290_ | \a[8] ) & ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))))))));
  assign new_n446_ = ((\a[5]  & ((new_n290_ & \a[8] ) | (~new_n290_ & ~\a[8] ) | ((~new_n291_ | ~\a[8] ) & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )))) & ((new_n290_ ^ \a[8] ) | (new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))) | (((\a[5]  & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )) & (~new_n292_ | (new_n291_ ^ \a[8] ))) | (~new_n349_ & (~\a[5]  | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )) | (new_n292_ & (~new_n291_ ^ \a[8] ))) & (\a[5]  | (~new_n292_ ^ (new_n291_ ^ \a[8] ))))) & (~\a[5]  | ((~new_n290_ | ~\a[8] ) & (new_n290_ | \a[8] ) & ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))) | ((~new_n290_ ^ \a[8] ) & (~new_n291_ | ~\a[8] ) & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )))) & (\a[5]  | ((new_n290_ ^ \a[8] ) ^ ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] ))))))) ^ (\a[5]  ^ ((~new_n289_ ^ ~\a[8] ) ^ ((new_n290_ & \a[8] ) | ((~new_n290_ | ~\a[8] ) & (new_n290_ | \a[8] ) & ((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )))))));
  assign new_n447_ = (\a[8]  ^ \a[11] ) ^ (new_n449_ ^ ((\a[5]  & (new_n278_ | (new_n44_ & \a[8] ) | (~new_n44_ & ~\a[8] )) & (~new_n278_ | (new_n44_ ^ \a[8] ))) | (~new_n448_ & (~\a[5]  | (~new_n278_ & (~new_n44_ | ~\a[8] ) & (new_n44_ | \a[8] )) | (new_n278_ & (~new_n44_ ^ \a[8] ))) & (\a[5]  | (~new_n278_ ^ (new_n44_ ^ \a[8] ))))));
  assign new_n448_ = (~new_n341_ | ~\a[5] ) & ((new_n341_ & \a[5] ) | (~new_n341_ & ~\a[5] ) | ((~new_n342_ | ~\a[5] ) & ((~new_n342_ & ~\a[5] ) | (new_n342_ & \a[5] ) | ((~new_n343_ | ~\a[5] ) & ((new_n343_ & \a[5] ) | (~new_n343_ & ~\a[5] ) | (~new_n344_ & (new_n345_ | ~new_n392_)))))));
  assign new_n449_ = (~new_n256_ | ~\a[14] ) & ((new_n256_ & \a[14] ) | (~new_n256_ & ~\a[14] ) | ((~new_n277_ | ~\a[14] ) & ((~new_n277_ & ~\a[14] ) | (new_n277_ & \a[14] ) | ((~new_n275_ | ~\a[14] ) & (new_n276_ | (~new_n275_ & ~\a[14] ) | (new_n275_ & \a[14] ))))));
  assign new_n450_ = ((~new_n340_ ^ \a[2] ) ^ ((new_n393_ & \a[2] ) | ((~new_n393_ | ~\a[2] ) & (new_n393_ | \a[2] ) & ((new_n394_ & \a[2] ) | ((~new_n394_ | ~\a[2] ) & (new_n394_ | \a[2] ) & ((\a[2]  & (new_n345_ | ~new_n392_) & (~new_n345_ | new_n392_)) | (~new_n395_ & (~\a[2]  | (~new_n345_ & new_n392_) | (new_n345_ & ~new_n392_)) & (\a[2]  | (~new_n345_ ^ new_n392_))))))))) & ((~new_n393_ ^ \a[2] ) ^ ((new_n394_ & \a[2] ) | ((~new_n394_ | ~\a[2] ) & (new_n394_ | \a[2] ) & ((\a[2]  & (new_n345_ | ~new_n392_) & (~new_n345_ | new_n392_)) | (~new_n395_ & (~\a[2]  | (~new_n345_ & new_n392_) | (new_n345_ & ~new_n392_)) & (\a[2]  | (~new_n345_ ^ new_n392_))))))) & ((~new_n394_ ^ \a[2] ) ^ ((\a[2]  & (new_n345_ | ~new_n392_) & (~new_n345_ | new_n392_)) | (~new_n395_ & (~\a[2]  | (~new_n345_ & new_n392_) | (new_n345_ & ~new_n392_)) & (\a[2]  | (~new_n345_ ^ new_n392_))))) & new_n451_ & (new_n395_ ^ (\a[2]  ^ (~new_n345_ ^ new_n392_)));
  assign new_n451_ = (((~new_n445_ | ~\a[2] ) & ((~new_n445_ & ~\a[2] ) | (new_n445_ & \a[2] ) | ((~new_n446_ | ~\a[2] ) & (new_n397_ | (new_n446_ & \a[2] ) | (~new_n446_ & ~\a[2] ))))) ^ (\a[2]  ^ (~new_n396_ ^ new_n347_))) & ((new_n445_ ^ ~\a[2] ) ^ ((new_n446_ & \a[2] ) | (~new_n397_ & (~new_n446_ | ~\a[2] ) & (new_n446_ | \a[2] )))) & new_n452_ & (new_n397_ ^ (new_n446_ ^ \a[2] ));
  assign new_n452_ = (~new_n454_ ^ (((new_n349_ | ~new_n401_) & (~new_n349_ | new_n401_) & \a[2] ) | (((new_n453_ & \a[2] ) | ((~new_n453_ | ~\a[2] ) & (new_n453_ | \a[2] ) & ((new_n402_ & \a[2] ) | (~new_n403_ & (~new_n402_ | ~\a[2] ) & (new_n402_ | \a[2] ))))) & ((~new_n349_ & new_n401_) | (new_n349_ & ~new_n401_) | ~\a[2] ) & ((~new_n349_ ^ new_n401_) | \a[2] )))) & (((~new_n453_ | ~\a[2] ) & ((new_n453_ & \a[2] ) | (~new_n453_ & ~\a[2] ) | ((~new_n402_ | ~\a[2] ) & (new_n403_ | (new_n402_ & \a[2] ) | (~new_n402_ & ~\a[2] ))))) ^ ((~new_n349_ ^ new_n401_) ^ \a[2] )) & ((~new_n453_ ^ \a[2] ) ^ ((new_n402_ & \a[2] ) | (~new_n403_ & (~new_n402_ | ~\a[2] ) & (new_n402_ | \a[2] )))) & (~new_n403_ | (new_n402_ ^ \a[2] )) & new_n455_ & (new_n403_ | (new_n402_ & \a[2] ) | (~new_n402_ & ~\a[2] ));
  assign new_n453_ = ~new_n399_ ^ (~new_n350_ ^ ~\a[5] );
  assign new_n454_ = \a[2]  ^ (((\a[5]  & (new_n292_ | (new_n291_ & \a[8] ) | (~new_n291_ & ~\a[8] )) & (~new_n292_ | (new_n291_ ^ \a[8] ))) | (~new_n349_ & (~\a[5]  | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] )) | (new_n292_ & (~new_n291_ ^ \a[8] ))) & (\a[5]  | (~new_n292_ ^ (new_n291_ ^ \a[8] ))))) ^ (\a[5]  ^ (((new_n291_ & \a[8] ) | (~new_n292_ & (~new_n291_ | ~\a[8] ) & (new_n291_ | \a[8] ))) ^ (~new_n290_ ^ ~\a[8] ))));
  assign new_n455_ = ((new_n456_ ^ \a[2] ) | (new_n457_ & \a[2] ) | ((new_n457_ | \a[2] ) & (~new_n457_ | ~\a[2] ) & ((new_n405_ & \a[2] ) | ((new_n405_ | \a[2] ) & (~new_n405_ | ~\a[2] ) & ((new_n483_ & \a[2] ) | (~new_n458_ & (~new_n483_ | ~\a[2] ) & (new_n483_ | \a[2] ))))))) & ((new_n456_ & \a[2] ) | (~new_n456_ & ~\a[2] ) | ((~new_n457_ | ~\a[2] ) & ((~new_n457_ & ~\a[2] ) | (new_n457_ & \a[2] ) | ((~new_n405_ | ~\a[2] ) & ((~new_n405_ & ~\a[2] ) | (new_n405_ & \a[2] ) | ((~new_n483_ | ~\a[2] ) & (new_n458_ | (new_n483_ & \a[2] ) | (~new_n483_ & ~\a[2] )))))))) & ((~new_n457_ ^ ~\a[2] ) | (new_n405_ & \a[2] ) | ((new_n405_ | \a[2] ) & (~new_n405_ | ~\a[2] ) & ((new_n483_ & \a[2] ) | (~new_n458_ & (~new_n483_ | ~\a[2] ) & (new_n483_ | \a[2] ))))) & ((~new_n457_ & ~\a[2] ) | (new_n457_ & \a[2] ) | ((~new_n405_ | ~\a[2] ) & ((~new_n405_ & ~\a[2] ) | (new_n405_ & \a[2] ) | ((~new_n483_ | ~\a[2] ) & (new_n458_ | (new_n483_ & \a[2] ) | (~new_n483_ & ~\a[2] )))))) & ((new_n405_ ^ ~\a[2] ) ^ ((new_n483_ & \a[2] ) | (~new_n458_ & (~new_n483_ | ~\a[2] ) & (new_n483_ | \a[2] )))) & (~new_n458_ | (new_n483_ ^ \a[2] )) & new_n460_ & (new_n458_ | (new_n483_ & \a[2] ) | (~new_n483_ & ~\a[2] ));
  assign new_n456_ = ~new_n351_ ^ new_n404_;
  assign new_n457_ = ~new_n400_ ^ (\a[5]  ^ (~new_n298_ ^ new_n352_));
  assign new_n458_ = (~\a[2]  | (~new_n459_ & new_n356_) | (new_n459_ & ~new_n356_)) & (((~new_n407_ | ~\a[2] ) & (((~new_n408_ | ~\a[2] ) & (new_n409_ | (~new_n408_ & ~\a[2] ) | (new_n408_ & \a[2] ))) | (~new_n407_ & ~\a[2] ) | (new_n407_ & \a[2] ))) | (\a[2]  & (new_n459_ | ~new_n356_) & (~new_n459_ | new_n356_)) | (~\a[2]  & (new_n459_ ^ new_n356_)));
  assign new_n459_ = ~new_n355_ ^ ~\a[5] ;
  assign new_n460_ = (((~new_n407_ | ~\a[2] ) & ((new_n407_ & \a[2] ) | (~new_n407_ & ~\a[2] ) | ((~new_n408_ | ~\a[2] ) & ((new_n408_ & \a[2] ) | (~new_n408_ & ~\a[2] ) | ((~new_n481_ | ~\a[2] ) & (new_n482_ | (new_n481_ & \a[2] ) | (~new_n481_ & ~\a[2] ))))))) ^ (\a[2]  ^ (new_n459_ ^ ~new_n356_))) & ((~new_n407_ ^ \a[2] ) ^ ((new_n408_ & \a[2] ) | ((~new_n408_ | ~\a[2] ) & (new_n408_ | \a[2] ) & ((new_n481_ & \a[2] ) | (~new_n482_ & (~new_n481_ | ~\a[2] ) & (new_n481_ | \a[2] )))))) & ((~new_n408_ ^ \a[2] ) ^ ((new_n481_ & \a[2] ) | (~new_n482_ & (~new_n481_ | ~\a[2] ) & (new_n481_ | \a[2] )))) & new_n461_ & (new_n482_ ^ (new_n481_ ^ \a[2] ));
  assign new_n461_ = ((new_n411_ ^ \a[2] ) | new_n412_ | (~new_n413_ & new_n444_)) & ((new_n411_ & \a[2] ) | (~new_n411_ & ~\a[2] ) | (~new_n412_ & (new_n413_ | ~new_n444_))) & (~new_n413_ | new_n444_) & (new_n413_ | ~new_n444_) & new_n462_ & (new_n479_ ^ new_n480_);
  assign new_n462_ = (~new_n463_ ^ (new_n417_ | (new_n441_ & ((new_n477_ & ~new_n421_) | (~new_n478_ & (new_n477_ | ~new_n421_) & (~new_n477_ | new_n421_)))))) & (~new_n441_ ^ ((new_n477_ & ~new_n421_) | (~new_n478_ & (new_n477_ | ~new_n421_) & (~new_n477_ | new_n421_)))) & (~new_n478_ | (~new_n477_ ^ new_n421_)) & new_n464_ & (new_n478_ | (~new_n477_ & new_n421_) | (new_n477_ & ~new_n421_));
  assign new_n463_ = ~new_n415_ ^ new_n443_;
  assign new_n464_ = ((~new_n423_ & (new_n425_ | ~new_n439_)) ^ (new_n422_ ^ ~new_n440_)) & (new_n425_ ^ new_n439_) & ~new_n475_ & new_n465_ & ~new_n476_;
  assign new_n465_ = (~new_n432_ | (~new_n430_ ^ new_n431_)) & new_n466_ & (new_n432_ | (~new_n430_ & new_n431_) | (new_n430_ & ~new_n431_));
  assign new_n466_ = (new_n467_ | (~new_n436_ & new_n437_) | (new_n438_ & (new_n436_ | ~new_n437_) & (~new_n436_ | new_n437_))) & (~new_n467_ | ((new_n436_ | ~new_n437_) & (~new_n438_ | (~new_n436_ & new_n437_) | (new_n436_ & ~new_n437_)))) & new_n468_ & (~new_n438_ | (~new_n436_ & new_n437_) | (new_n436_ & ~new_n437_)) & ~new_n474_ & (new_n438_ | (~new_n436_ ^ new_n437_));
  assign new_n467_ = new_n435_ ^ (~\a[2]  ^ (new_n434_ & (~new_n60_ | ~new_n433_)));
  assign new_n468_ = (~new_n469_ | ~new_n470_ | ~new_n471_) & \a[0]  & \b[0]  & (~new_n472_ | ~new_n473_);
  assign new_n469_ = ~\a[5]  & ~\a[6]  & ~\a[7]  & ~\a[8]  & ~\a[1]  & ~\a[2]  & ~\a[3]  & ~\a[4] ;
  assign new_n470_ = ~\a[11]  & ~\a[12]  & ~\a[15]  & ~\a[16]  & ~\a[9]  & ~\a[10]  & ~\a[13]  & ~\a[14] ;
  assign new_n471_ = ~\a[21]  & ~\a[22]  & ~\a[23]  & ~\a[24]  & ~\a[17]  & ~\a[18]  & ~\a[19]  & ~\a[20] ;
  assign new_n472_ = ~\b[1]  & ~\b[2]  & ~\b[3]  & ~\b[4] ;
  assign new_n473_ = ~\b[9]  & ~\b[10]  & ~\b[11]  & ~\b[12]  & ~\b[5]  & ~\b[6]  & ~\b[7]  & ~\b[8] ;
  assign new_n474_ = ((\b[2]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[1]  & ~\a[0]  & \a[1] ) | (\b[0]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | ((~\b[2]  ^ (\b[0]  | ~\b[1] )) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[0]  & ~\a[0]  & \a[1] ) | (\b[1]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | ((\b[0]  ^ \b[1] ) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | ~\a[2]  | (\a[0]  & \b[0] )) & ((\b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (~\a[2]  ^ ((~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] ) & (((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))))) | ((~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\a[2]  | (\b[1]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[3]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[2]  & ~\a[0]  & \a[1] ) | (((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )) & ((\b[2]  ^ \b[3] ) | (\b[1]  & (\b[0]  | \b[2] ))) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] ))) & (\a[2]  | ((~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] ) & (((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))))) | (\a[2]  & (~\a[0]  | ~\b[0]  | ((~\b[1]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & ((~\b[0]  ^ \b[1] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))))) | (((~\b[2]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[1]  | \a[0]  | ~\a[1] ) & (~\b[0]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & ((\b[2]  ^ (\b[0]  | ~\b[1] )) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))) ? ((\b[0]  & ~\a[0]  & \a[1] ) | (\b[1]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | ((\b[0]  ^ \b[1] ) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] ))) : ~\a[2] ));
  assign new_n475_ = (~new_n427_ ^ (~new_n377_ ^ new_n426_)) ^ ((~new_n428_ & new_n429_) | ((new_n428_ | ~new_n429_) & (~new_n428_ | new_n429_) & ((~new_n430_ & new_n431_) | (~new_n432_ & (new_n430_ | ~new_n431_) & (~new_n430_ | new_n431_)))));
  assign new_n476_ = (~new_n428_ ^ new_n429_) ^ ((~new_n430_ & new_n431_) | (~new_n432_ & (new_n430_ | ~new_n431_) & (~new_n430_ | new_n431_)));
  assign new_n477_ = ~new_n369_ ^ new_n420_;
  assign new_n478_ = (~new_n422_ | new_n440_) & ((~new_n423_ & (new_n425_ | ~new_n439_)) | (new_n422_ & ~new_n440_) | (~new_n422_ & new_n440_));
  assign new_n479_ = (~new_n415_ | new_n443_) & ((~new_n417_ & (new_n419_ | ~new_n441_)) | (new_n415_ & ~new_n443_) | (~new_n415_ & new_n443_));
  assign new_n480_ = ~new_n442_ ^ (~new_n363_ ^ new_n414_);
  assign new_n481_ = ~new_n358_ ^ new_n410_;
  assign new_n482_ = (~new_n411_ | ~\a[2] ) & ((new_n411_ & \a[2] ) | (~new_n411_ & ~\a[2] ) | (~new_n412_ & (new_n413_ | ~new_n444_)));
  assign new_n483_ = (new_n354_ ^ \a[5] ) ^ ((new_n355_ & \a[5] ) | (~new_n356_ & (~new_n355_ | ~\a[5] ) & (new_n355_ | \a[5] )));
  assign new_n484_ = \a[5]  ^ (~new_n278_ ^ (new_n44_ ^ \a[8] ));
endmodule


