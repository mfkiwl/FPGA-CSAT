// Benchmark "multiplier_907_sat" written by ABC on Fri Jan 27 15:09:01 2023

module multiplier_907_sat ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    sat  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ;
  output sat;
  wire new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_, new_n24_,
    new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_, new_n31_,
    new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_, new_n38_,
    new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_, new_n45_,
    new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_, new_n52_,
    new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_, new_n59_,
    new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_,
    new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n73_,
    new_n74_;
  assign sat = ~new_n18_ & new_n60_ & (~new_n43_ ^ (~new_n57_ ^ (~new_n58_ ^ (\a[2]  ^ \a[5] ))));
  assign new_n18_ = (new_n41_ ^ \a[5] ) ^ ((~new_n19_ & new_n40_) | (new_n37_ & \a[5] ));
  assign new_n19_ = (~new_n33_ | ~\a[5] ) & (((new_n32_ | ~new_n36_) & ((~new_n28_ & (new_n20_ | ~new_n31_)) | (~new_n32_ & new_n36_) | (new_n32_ & ~new_n36_))) | (new_n33_ & \a[5] ) | (~new_n33_ & ~\a[5] ));
  assign new_n20_ = (~new_n24_ | (\a[5]  ^ (new_n23_ & (~new_n21_ | ~new_n22_)))) & ((~new_n25_ & (new_n26_ | ~new_n27_)) | (new_n24_ & (~\a[5]  ^ (new_n23_ & (~new_n21_ | ~new_n22_)))) | (~new_n24_ & (~\a[5]  | ~new_n23_ | (new_n21_ & new_n22_)) & (\a[5]  | (new_n23_ & (~new_n21_ | ~new_n22_)))));
  assign new_n21_ = (~\a[2]  | ~\a[3] ) & (\a[2]  | \a[3] ) & (\a[4]  | \a[5] ) & (~\a[4]  | ~\a[5] );
  assign new_n22_ = (\b[3]  ^ \b[4] ) ^ ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] )));
  assign new_n23_ = (~\b[2]  | (~\a[3]  ^ ~\a[4] ) | (\a[2]  ^ \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )) & (~\b[3]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[4]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] ));
  assign new_n24_ = ((\b[0]  & (~\a[5]  ^ \a[6] ) & (\a[6]  | \a[7] ) & (~\a[6]  | ~\a[7] )) | (\b[1]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  ^ ~\a[8] )) | ((~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] ) & (\b[0]  ^ \b[1] ))) ^ (\a[8]  & \b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ));
  assign new_n25_ = \b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (~\b[0]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\b[0]  ^ \b[1] ) | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )) & \a[5]  & (~\b[0]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] )) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (\a[2]  ^ \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )) & ((\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | ((\b[0]  | ~\b[1] ) ^ \b[2] )) & (~\b[2]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[1]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ));
  assign new_n26_ = \a[5]  ^ (((\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (~\a[3]  ^ ~\a[4] ) | (\a[2]  ^ \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )) & (~\b[3]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[2]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )));
  assign new_n27_ = (\b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] )) ^ ((~\b[0]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\b[0]  ^ \b[1] ) | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )) & \a[5]  & (~\b[0]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] )) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (\a[2]  ^ \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )) & ((\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | ((\b[0]  | ~\b[1] ) ^ \b[2] )) & (~\b[2]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[1]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )));
  assign new_n28_ = new_n30_ & (~\a[5]  ^ (((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~new_n29_ ^ ~\b[4] )) & (~\b[3]  | (\a[3]  ^ \a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )) & (~\b[4]  | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] ) | (~\a[2]  ^ ~\a[3] ))));
  assign new_n29_ = (~\b[3]  | ~\b[4] ) & ((\b[3]  & \b[4] ) | (~\b[3]  & ~\b[4] ) | ((~\b[2]  | ~\b[3] ) & ((~\b[2]  & ~\b[3] ) | (\b[2]  & \b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] ))));
  assign new_n30_ = ((~\b[0]  | (\a[5]  ^ \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[6]  ^ ~\a[7] )) & (~\b[1]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[2]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))) ^ (~\a[8]  | ((~\b[0]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\b[0]  ^ \b[1] )) & \a[8]  & (~\b[0]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ))));
  assign new_n31_ = new_n30_ ^ (~\a[5]  ^ (((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~new_n29_ ^ ~\b[4] )) & (~\b[3]  | (\a[3]  ^ \a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )) & (~\b[4]  | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] ) | (~\a[2]  ^ ~\a[3] ))));
  assign new_n32_ = \a[5]  ^ (~\b[4]  | ((new_n29_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] ))));
  assign new_n33_ = ~new_n34_ ^ ((\a[8]  & ~\b[1] ) ^ (~new_n35_ | (new_n22_ & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] ))));
  assign new_n34_ = (~\a[8]  | ~\b[0]  | (\b[0]  & (~\a[5]  ^ \a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] ) & (\a[6]  ^ ~\a[7] )) | (\b[1]  & (~\a[5]  ^ \a[6] ) & (\a[6]  | \a[7] ) & (~\a[6]  | ~\a[7] )) | (\b[2]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  ^ ~\a[8] )) | ((~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] ) & (~\b[2]  ^ (\b[0]  | ~\b[1] ))) | (\b[0]  & (~\a[5]  ^ \a[6] ) & (\a[6]  | \a[7] ) & (~\a[6]  | ~\a[7] )) | (\b[1]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  ^ ~\a[8] )) | ((~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] ) & (\b[0]  ^ \b[1] )) | (\b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ))) & ((\a[8]  ^ (((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[2]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (\a[5]  ^ \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[6]  ^ ~\a[7] )))) | (\a[8]  & \b[0]  & (~\b[0]  | (\a[5]  ^ \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[6]  ^ ~\a[7] )) & (~\b[1]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[2]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\b[0]  ^ \b[1] )) & (~\b[0]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ))) | ((~\a[8]  | ~\b[0] ) & ((\b[0]  & (~\a[5]  ^ \a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] ) & (\a[6]  ^ ~\a[7] )) | (\b[1]  & (~\a[5]  ^ \a[6] ) & (\a[6]  | \a[7] ) & (~\a[6]  | ~\a[7] )) | (\b[2]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  ^ ~\a[8] )) | ((~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] ) & (~\b[2]  ^ (\b[0]  | ~\b[1] ))) | (\b[0]  & (~\a[5]  ^ \a[6] ) & (\a[6]  | \a[7] ) & (~\a[6]  | ~\a[7] )) | (\b[1]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  ^ ~\a[8] )) | ((~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] ) & (\b[0]  ^ \b[1] )) | ~\a[8]  | (\b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] )))));
  assign new_n35_ = (~\b[3]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[4]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[2]  | (\a[5]  ^ \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[6]  ^ ~\a[7] ));
  assign new_n36_ = (~\a[8]  ^ (((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[2]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (\a[5]  ^ \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[6]  ^ ~\a[7] )))) ^ ((\a[8]  & \b[0] ) ^ ((~\b[0]  | (\a[5]  ^ \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[6]  ^ ~\a[7] )) & (~\b[1]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[2]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\b[0]  ^ \b[1] )) & \a[8]  & (~\b[0]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ))));
  assign new_n37_ = ~new_n39_ ^ (~new_n38_ ^ (\a[8]  & ~\b[2] ));
  assign new_n38_ = ((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~new_n29_ ^ ~\b[4] )) & (~\b[3]  | (~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[6]  ^ ~\a[7] )) & (~\b[4]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] ));
  assign new_n39_ = (new_n34_ | (\a[8]  & ~\b[1]  & (~new_n35_ | (new_n22_ & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] )))) | ((~\a[8]  | \b[1] ) & new_n35_ & (~new_n22_ | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )))) & (~\a[8]  | ~\b[1]  | ~new_n35_ | (new_n22_ & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] )));
  assign new_n40_ = \a[5]  ^ (~new_n39_ ^ (~new_n38_ ^ (\a[8]  & ~\b[2] )));
  assign new_n41_ = new_n42_ ^ ((new_n39_ | (~new_n38_ & \a[8]  & ~\b[2] ) | (new_n38_ & (~\a[8]  | \b[2] ))) & (~new_n38_ | ~\a[8]  | ~\b[2] ));
  assign new_n42_ = (\a[8]  & ~\b[3] ) ^ (~\b[4]  | ((new_n29_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[6]  ^ ~\a[7] ))));
  assign new_n43_ = (~\a[2]  | (~new_n46_ & (new_n19_ ^ (new_n37_ ^ \a[5] )) & ~new_n44_ & ~new_n55_)) & (((~new_n41_ | ~\a[5] ) & (new_n41_ | \a[5] ) & ((new_n37_ & \a[5] ) | (~new_n19_ & (~new_n37_ | ~\a[5] ) & (new_n37_ | \a[5] )))) | ((~new_n41_ ^ \a[5] ) & (~new_n37_ | ~\a[5] ) & (new_n19_ | (new_n37_ & \a[5] ) | (~new_n37_ & ~\a[5] ))) | (~\a[2]  & (~new_n46_ | ~new_n55_ | (~new_n19_ & (~new_n37_ | ~\a[5] ) & (new_n37_ | \a[5] )) | (new_n19_ & (~new_n37_ ^ \a[5] )))));
  assign new_n44_ = new_n45_ ^ (new_n28_ | (~new_n20_ & new_n31_));
  assign new_n45_ = new_n36_ ^ (~\a[5]  ^ (~\b[4]  | (((\a[3]  ^ \a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )) & (new_n29_ | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )))));
  assign new_n46_ = ((\a[2]  & (new_n20_ | ~new_n31_) & (~new_n20_ | new_n31_)) | (((new_n47_ & \a[2] ) | (~new_n48_ & (~new_n47_ | ~\a[2] ) & (new_n47_ | \a[2] ))) & (~\a[2]  | (~new_n20_ & new_n31_) | (new_n20_ & ~new_n31_)) & (\a[2]  | (~new_n20_ ^ new_n31_)))) & (~\a[2]  ^ (~new_n45_ ^ (new_n28_ | (~new_n20_ & new_n31_))));
  assign new_n47_ = (new_n25_ | (~new_n26_ & new_n27_)) ^ (new_n24_ ^ (~\a[5]  ^ (new_n23_ & (~new_n21_ | ~new_n22_))));
  assign new_n48_ = (new_n49_ | (~new_n26_ & new_n27_) | (new_n26_ & ~new_n27_)) & (((new_n50_ | ~new_n51_) & (((new_n52_ | ~new_n53_) & ((~new_n52_ & new_n53_) | (new_n52_ & ~new_n53_) | ~new_n54_)) | (new_n50_ & ~new_n51_) | (~new_n50_ & new_n51_))) | (~new_n49_ & (new_n26_ | ~new_n27_) & (~new_n26_ | new_n27_)) | (new_n49_ & (new_n26_ ^ new_n27_)));
  assign new_n49_ = \a[2]  ^ (~\b[4]  | ((((~\b[3]  | ~\b[4] ) & ((\b[3]  & \b[4] ) | (~\b[3]  & ~\b[4] ) | ((~\b[2]  | ~\b[3] ) & ((~\b[2]  & ~\b[3] ) | (\b[2]  & \b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] ))))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (\a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))));
  assign new_n50_ = \a[2]  ^ ((~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | (~\b[4]  ^ ((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))))) & (~\b[3]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[4]  | \a[0]  | ~\a[1] ));
  assign new_n51_ = (~\a[5]  | ((~\b[0]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\b[0]  ^ \b[1] )) & \a[5]  & (~\b[0]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] )))) ^ ((~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (\a[2]  ^ \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )) & (~\b[1]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[2]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n52_ = \a[2]  ^ ((~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] )))) | ((~\b[3]  ^ \b[4] ) & (~\b[2]  | ~\b[3] ) & ((~\b[2]  & ~\b[3] ) | (\b[2]  & \b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[4]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[3]  | \a[0]  | ~\a[1] ));
  assign new_n53_ = ((\b[0]  & (~\a[2]  ^ \a[3] ) & (\a[3]  | \a[4] ) & (~\a[3]  | ~\a[4] )) | (\b[1]  & (~\a[2]  | ~\a[3] ) & (\a[2]  | \a[3] ) & (\a[4]  ^ ~\a[5] )) | ((~\a[2]  | ~\a[3] ) & (\a[2]  | \a[3] ) & (\a[4]  | \a[5] ) & (~\a[4]  | ~\a[5] ) & (\b[0]  ^ \b[1] ))) ^ (\a[5]  & \b[0]  & (~\a[2]  | ~\a[3] ) & (\a[2]  | \a[3] ));
  assign new_n54_ = ((\b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] )) | (\a[2]  & (~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] ) & (((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))) | (~\a[2]  & ((\b[1]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[3]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[2]  & ~\a[0]  & \a[1] ) | (((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )) & ((\b[2]  ^ \b[3] ) | (\b[1]  & (\b[0]  | \b[2] ))) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] ))))) & ((\b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (~\a[2]  ^ ((~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] ) & (((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))))) | ((~\b[1]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & ((~\b[0]  ^ \b[1] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[0]  | \a[0]  | ~\a[1] ) & (~\b[2]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[1]  | \a[0]  | ~\a[1] ) & (~\b[0]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & ((\b[2]  ^ (\b[0]  | ~\b[1] )) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & \a[2]  & (~\a[0]  | ~\b[0] )));
  assign new_n55_ = new_n56_ ^ ((~new_n32_ & new_n36_) | ((new_n28_ | (~new_n20_ & new_n31_)) & (new_n32_ | ~new_n36_) & (~new_n32_ | new_n36_)));
  assign new_n56_ = \a[5]  ^ (~new_n34_ ^ ((\a[8]  & ~\b[1] ) ^ (~new_n35_ | (new_n22_ & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] )))));
  assign new_n57_ = (~\a[8]  | \b[4] ) ^ ((~new_n41_ | ~\a[5] ) & ((new_n41_ & \a[5] ) | (~new_n41_ & ~\a[5] ) | ((new_n19_ | ~new_n40_) & (~new_n37_ | ~\a[5] ))));
  assign new_n58_ = (new_n59_ | ((\a[8]  & ~\b[3] ) ^ (~\b[4]  | (((~\a[5]  ^ ~\a[6] ) | (\a[6]  ^ \a[7] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )) & (new_n29_ | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )))))) & (~\a[8]  | ~\b[3]  | (\b[4]  & (((\a[5]  ^ ~\a[6] ) & (~\a[6]  ^ \a[7] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] )) | (~new_n29_ & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] )))));
  assign new_n59_ = (new_n39_ | (~new_n38_ & \a[8]  & ~\b[2] ) | (new_n38_ & (~\a[8]  | \b[2] ))) & (~new_n38_ | ~\a[8]  | ~\b[2] );
  assign new_n60_ = new_n74_ & ~new_n62_ & ~new_n61_ & new_n63_ & ~new_n73_ & (new_n19_ ^ new_n40_);
  assign new_n61_ = ((new_n47_ & \a[2] ) | (~new_n48_ & (~new_n47_ | ~\a[2] ) & (new_n47_ | \a[2] ))) & (~\a[2]  | (~new_n20_ & new_n31_) | (new_n20_ & ~new_n31_)) & (\a[2]  | (~new_n20_ ^ new_n31_));
  assign new_n62_ = (~new_n47_ | ~\a[2] ) & (new_n48_ | (new_n47_ & \a[2] ) | (~new_n47_ & ~\a[2] )) & (~\a[2]  ^ (~new_n20_ ^ new_n31_));
  assign new_n63_ = (~new_n48_ | (~new_n47_ ^ ~\a[2] )) & (new_n48_ | (~new_n47_ & ~\a[2] ) | (new_n47_ & \a[2] )) & ~new_n64_ & ~new_n65_ & ~new_n66_ & new_n67_;
  assign new_n64_ = ((~new_n50_ & new_n51_) | (((~new_n52_ & new_n53_) | ((new_n52_ | ~new_n53_) & (~new_n52_ | new_n53_) & new_n54_)) & (~new_n50_ | new_n51_) & (new_n50_ | ~new_n51_))) ^ (~new_n49_ ^ (~new_n26_ ^ new_n27_));
  assign new_n65_ = (~new_n50_ ^ new_n51_) ^ ((~new_n52_ & new_n53_) | (new_n54_ & (~new_n52_ | new_n53_) & (new_n52_ | ~new_n53_)));
  assign new_n66_ = new_n54_ ^ (~new_n52_ ^ new_n53_);
  assign new_n67_ = (new_n68_ | ~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~new_n68_ | (\b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ))) & ~new_n69_ & ~new_n70_ & ~new_n71_ & new_n72_;
  assign new_n68_ = \a[2]  ^ ((~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((\b[2]  ^ ~\b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] ) & (~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )));
  assign new_n69_ = \a[2]  ? ((\b[1]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | ((~\b[0]  ^ ~\b[1] ) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[0]  & ~\a[0]  & \a[1] )) : ((\b[2]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[1]  & ~\a[0]  & \a[1] ) | (\b[0]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] ) & (~\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n70_ = (~\b[2]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[1]  | \a[0]  | ~\a[1] ) & (~\b[0]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[1]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & ((\b[0]  ^ ~\b[1] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[0]  | \a[0]  | ~\a[1] );
  assign new_n71_ = ~\a[7]  & ~\a[8]  & ~\a[5]  & ~\a[6]  & ~\a[1]  & ~\a[2]  & ~\a[3]  & ~\a[4] ;
  assign new_n72_ = \a[0]  & \b[0]  & (\b[2]  | \b[3]  | \b[1]  | \b[4] );
  assign new_n73_ = (~new_n56_ ^ ((~new_n32_ & new_n36_) | ((new_n28_ | (~new_n20_ & new_n31_)) & (new_n32_ | ~new_n36_) & (~new_n32_ | new_n36_)))) ^ (~\a[2]  | ((new_n28_ | (~new_n20_ & new_n31_)) ^ (~new_n32_ ^ new_n36_)));
  assign new_n74_ = ((\a[2]  & (new_n20_ | ~new_n31_) & (~new_n20_ | new_n31_)) | (((new_n47_ & \a[2] ) | (~new_n48_ & (~new_n47_ | ~\a[2] ) & (new_n47_ | \a[2] ))) & (~\a[2]  | (~new_n20_ & new_n31_) | (new_n20_ & ~new_n31_)) & (\a[2]  | (~new_n20_ ^ new_n31_)))) ^ (~\a[2]  ^ (~new_n45_ ^ (new_n28_ | (~new_n20_ & new_n31_))));
endmodule


