// Benchmark "multiplier_7485671_sat" written by ABC on Fri Nov 11 15:27:54 2022

module multiplier_7485671_sat ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \b[0] , \b[1] , \b[2] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] ,
    \b[11] ,
    sat  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \b[0] , \b[1] ,
    \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] ;
  output sat;
  wire new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_,
    new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_,
    new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_;
  assign sat = (new_n357_ ^ ((~new_n38_ | ~\a[2] ) & ((new_n38_ & \a[2] ) | (~new_n38_ & ~\a[2] ) | ((~new_n398_ | ~\a[2] ) & (((~new_n399_ | ~\a[2] ) & ((new_n399_ & \a[2] ) | (~new_n399_ & ~\a[2] ) | ((~new_n400_ | ~\a[2] ) & (new_n309_ | (new_n400_ & \a[2] ) | (~new_n400_ & ~\a[2] ))))) | (new_n398_ & \a[2] ) | (~new_n398_ & ~\a[2] )))))) & ((~new_n38_ ^ \a[2] ) ^ ((new_n398_ & \a[2] ) | (((new_n399_ & \a[2] ) | ((~new_n399_ | ~\a[2] ) & (new_n399_ | \a[2] ) & ((new_n400_ & \a[2] ) | (~new_n309_ & (~new_n400_ | ~\a[2] ) & (new_n400_ | \a[2] ))))) & (~new_n398_ | ~\a[2] ) & (new_n398_ | \a[2] )))) & (((~new_n399_ | ~\a[2] ) & ((new_n399_ & \a[2] ) | (~new_n399_ & ~\a[2] ) | ((~new_n400_ | ~\a[2] ) & (new_n309_ | (new_n400_ & \a[2] ) | (~new_n400_ & ~\a[2] ))))) ^ (new_n398_ ^ \a[2] )) & ((~new_n399_ ^ \a[2] ) ^ ((new_n400_ & \a[2] ) | (~new_n309_ & (~new_n400_ | ~\a[2] ) & (new_n400_ | \a[2] )))) & new_n366_ & (new_n309_ ^ (new_n400_ ^ \a[2] ));
  assign new_n38_ = ~new_n39_ ^ (~new_n302_ ^ ~\a[5] );
  assign new_n39_ = (~\a[5]  | (~new_n40_ & new_n242_) | (new_n40_ & ~new_n242_)) & (((~new_n250_ | ~\a[5] ) & ((new_n250_ & \a[5] ) | (~new_n250_ & ~\a[5] ) | ((~new_n251_ | ~\a[5] ) & (((~new_n253_ | ~\a[5] ) & (new_n254_ | (new_n253_ & \a[5] ) | (~new_n253_ & ~\a[5] ))) | (new_n251_ & \a[5] ) | (~new_n251_ & ~\a[5] ))))) | (\a[5]  & (new_n40_ | ~new_n242_) & (~new_n40_ | new_n242_)) | (~\a[5]  & (new_n40_ ^ new_n242_)));
  assign new_n40_ = (~\a[8]  | ((~new_n178_ | ~\a[11] ) & (new_n178_ | \a[11] ) & ((new_n241_ & \a[11] ) | (~new_n41_ & (~new_n241_ | ~\a[11] ) & (new_n241_ | \a[11] )))) | ((~new_n178_ ^ \a[11] ) & (~new_n241_ | ~\a[11] ) & (new_n41_ | (new_n241_ & \a[11] ) | (~new_n241_ & ~\a[11] )))) & (((~\a[8]  | (~new_n41_ & (~new_n241_ | ~\a[11] ) & (new_n241_ | \a[11] )) | (new_n41_ & (~new_n241_ ^ \a[11] ))) & (((~new_n195_ | ~\a[8] ) & ((new_n195_ & \a[8] ) | (~new_n195_ & ~\a[8] ) | ((~new_n196_ | ~\a[8] ) & (new_n199_ | (new_n196_ & \a[8] ) | (~new_n196_ & ~\a[8] ))))) | (\a[8]  & (new_n41_ | (new_n241_ & \a[11] ) | (~new_n241_ & ~\a[11] )) & (~new_n41_ | (new_n241_ ^ \a[11] ))) | (~\a[8]  & (new_n41_ ^ (new_n241_ ^ \a[11] ))))) | (\a[8]  & ((new_n178_ & \a[11] ) | (~new_n178_ & ~\a[11] ) | ((~new_n241_ | ~\a[11] ) & (new_n41_ | (new_n241_ & \a[11] ) | (~new_n241_ & ~\a[11] )))) & ((new_n178_ ^ \a[11] ) | (new_n241_ & \a[11] ) | (~new_n41_ & (~new_n241_ | ~\a[11] ) & (new_n241_ | \a[11] )))) | (~\a[8]  & ((~new_n178_ ^ \a[11] ) ^ ((new_n241_ & \a[11] ) | (~new_n41_ & (~new_n241_ | ~\a[11] ) & (new_n241_ | \a[11] ))))));
  assign new_n41_ = (~\a[11]  | ((~new_n151_ | ~\a[14] ) & (new_n151_ | \a[14] ) & ((new_n174_ & \a[14] ) | (((\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~new_n175_ & (~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (\a[14]  | (~new_n163_ ^ new_n177_)))) & (~new_n174_ | ~\a[14] ) & (new_n174_ | \a[14] )))) | ((~new_n151_ ^ \a[14] ) & (~new_n174_ | ~\a[14] ) & (((~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (new_n175_ | (\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~\a[14]  & (new_n163_ ^ new_n177_)))) | (new_n174_ & \a[14] ) | (~new_n174_ & ~\a[14] )))) & (((~\a[11]  | (((\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~new_n175_ & (~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (\a[14]  | (~new_n163_ ^ new_n177_)))) & (~new_n174_ | ~\a[14] ) & (new_n174_ | \a[14] )) | ((~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (new_n175_ | (\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~\a[14]  & (new_n163_ ^ new_n177_))) & (~new_n174_ ^ \a[14] ))) & (((~\a[11]  | (~new_n175_ & (~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (\a[14]  | (~new_n163_ ^ new_n177_))) | (new_n175_ & (~\a[14]  ^ (~new_n163_ ^ new_n177_)))) & (new_n42_ | (\a[11]  & (new_n175_ | (\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~\a[14]  & (new_n163_ ^ new_n177_))) & (~new_n175_ | (\a[14]  ^ (~new_n163_ ^ new_n177_)))) | (~\a[11]  & (new_n175_ ^ (\a[14]  ^ (~new_n163_ ^ new_n177_)))))) | (\a[11]  & (((~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (new_n175_ | (\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~\a[14]  & (new_n163_ ^ new_n177_)))) | (new_n174_ & \a[14] ) | (~new_n174_ & ~\a[14] )) & ((\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~new_n175_ & (~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (\a[14]  | (~new_n163_ ^ new_n177_))) | (new_n174_ ^ \a[14] ))) | (~\a[11]  & (((~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (new_n175_ | (\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~\a[14]  & (new_n163_ ^ new_n177_)))) ^ (new_n174_ ^ \a[14] ))))) | (\a[11]  & ((new_n151_ & \a[14] ) | (~new_n151_ & ~\a[14] ) | ((~new_n174_ | ~\a[14] ) & (((~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (new_n175_ | (\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~\a[14]  & (new_n163_ ^ new_n177_)))) | (new_n174_ & \a[14] ) | (~new_n174_ & ~\a[14] )))) & ((new_n151_ ^ \a[14] ) | (new_n174_ & \a[14] ) | (((\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~new_n175_ & (~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (\a[14]  | (~new_n163_ ^ new_n177_)))) & (~new_n174_ | ~\a[14] ) & (new_n174_ | \a[14] )))) | (~\a[11]  & ((~new_n151_ ^ \a[14] ) ^ ((new_n174_ & \a[14] ) | (((\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~new_n175_ & (~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (\a[14]  | (~new_n163_ ^ new_n177_)))) & (~new_n174_ | ~\a[14] ) & (new_n174_ | \a[14] ))))));
  assign new_n42_ = (~\a[11]  | (new_n123_ & (new_n143_ | (new_n149_ & ((new_n145_ & ~new_n150_) | (~new_n146_ & (~new_n145_ | new_n150_) & (new_n145_ | ~new_n150_)))))) | (~new_n123_ & ~new_n143_ & (~new_n149_ | ((~new_n145_ | new_n150_) & (new_n146_ | (new_n145_ & ~new_n150_) | (~new_n145_ & new_n150_)))))) & (((~\a[11]  | (new_n149_ & ((new_n145_ & ~new_n150_) | (~new_n146_ & (~new_n145_ | new_n150_) & (new_n145_ | ~new_n150_)))) | (~new_n149_ & (~new_n145_ | new_n150_) & (new_n146_ | (new_n145_ & ~new_n150_) | (~new_n145_ & new_n150_)))) & (((~\a[11]  | (~new_n146_ & (~new_n145_ | new_n150_) & (new_n145_ | ~new_n150_)) | (new_n146_ & (~new_n145_ ^ ~new_n150_))) & (new_n43_ | (\a[11]  & (new_n146_ | (new_n145_ & ~new_n150_) | (~new_n145_ & new_n150_)) & (~new_n146_ | (new_n145_ ^ ~new_n150_))) | (~\a[11]  & (new_n146_ ^ (new_n145_ ^ ~new_n150_))))) | (\a[11]  & (~new_n149_ | ((~new_n145_ | new_n150_) & (new_n146_ | (new_n145_ & ~new_n150_) | (~new_n145_ & new_n150_)))) & (new_n149_ | (new_n145_ & ~new_n150_) | (~new_n146_ & (~new_n145_ | new_n150_) & (new_n145_ | ~new_n150_)))) | (~\a[11]  & (~new_n149_ ^ ((new_n145_ & ~new_n150_) | (~new_n146_ & (~new_n145_ | new_n150_) & (new_n145_ | ~new_n150_))))))) | (\a[11]  & (~new_n123_ | (~new_n143_ & (~new_n149_ | ((~new_n145_ | new_n150_) & (new_n146_ | (new_n145_ & ~new_n150_) | (~new_n145_ & new_n150_)))))) & (new_n123_ | new_n143_ | (new_n149_ & ((new_n145_ & ~new_n150_) | (~new_n146_ & (~new_n145_ | new_n150_) & (new_n145_ | ~new_n150_)))))) | (~\a[11]  & (~new_n123_ ^ (new_n143_ | (new_n149_ & ((new_n145_ & ~new_n150_) | (~new_n146_ & (~new_n145_ | new_n150_) & (new_n145_ | ~new_n150_))))))));
  assign new_n43_ = (~new_n44_ | new_n122_) & ((~new_n90_ & (~new_n121_ | (~new_n93_ & (new_n97_ | ~new_n120_)))) | (new_n44_ & ~new_n122_) | (~new_n44_ & new_n122_));
  assign new_n44_ = new_n80_ ^ (new_n45_ | (new_n79_ & ((~new_n89_ & (new_n53_ | (~new_n51_ & new_n63_) | (new_n51_ & ~new_n63_)) & (~new_n53_ | (~new_n51_ ^ new_n63_))) | (~new_n64_ & (new_n89_ | (~new_n53_ & (new_n51_ | ~new_n63_) & (~new_n51_ | new_n63_)) | (new_n53_ & (new_n51_ ^ new_n63_))) & (~new_n89_ | (~new_n53_ ^ (~new_n51_ ^ new_n63_)))))));
  assign new_n45_ = ~new_n61_ & ((~new_n46_ & new_n49_) | (new_n46_ & ~new_n49_) | ((new_n51_ | ~new_n63_) & (new_n53_ | (~new_n51_ & new_n63_) | (new_n51_ & ~new_n63_)))) & ((~new_n46_ ^ new_n49_) | (~new_n51_ & new_n63_) | (~new_n53_ & (new_n51_ | ~new_n63_) & (~new_n51_ | new_n63_)));
  assign new_n46_ = ~new_n47_ ^ new_n48_;
  assign new_n47_ = \a[20]  ^ (((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[2]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[3]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )));
  assign new_n48_ = (\b[0]  & (\a[20]  ^ \a[21] )) ^ ((~\b[0]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[1]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[20]  & (~\b[0]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[0]  | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[1]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[2]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n49_ = \a[17]  ^ ((~new_n50_ | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )) & (~\b[4]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & (~\b[5]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[6]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  ^ \a[17] )));
  assign new_n50_ = (\b[5]  ^ \b[6] ) ^ ((\b[4]  & \b[5] ) | (((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))) & (~\b[4]  | ~\b[5] ) & (\b[4]  | \b[5] )));
  assign new_n51_ = \a[17]  ^ ((~new_n52_ | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )) & (~\b[3]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & (~\b[4]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[5]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  ^ \a[17] )));
  assign new_n52_ = ((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))) ^ (\b[4]  ^ \b[5] );
  assign new_n53_ = (~new_n57_ | (\a[17]  ^ (new_n56_ & (~new_n54_ | ~new_n55_)))) & ((~new_n58_ & (new_n59_ | ~new_n60_)) | (new_n57_ & (~\a[17]  ^ (new_n56_ & (~new_n54_ | ~new_n55_)))) | (~new_n57_ & (~\a[17]  | ~new_n56_ | (new_n54_ & new_n55_)) & (\a[17]  | (new_n56_ & (~new_n54_ | ~new_n55_)))));
  assign new_n54_ = (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ) & (\a[16]  | \a[17] ) & (~\a[16]  | ~\a[17] );
  assign new_n55_ = (\b[3]  ^ \b[4] ) ^ ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] )));
  assign new_n56_ = (~\b[2]  | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[3]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[4]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] ));
  assign new_n57_ = ((\b[0]  & (\a[18]  | \a[19] ) & (~\a[18]  | ~\a[19] ) & (\a[17]  ^ ~\a[18] )) | (\b[1]  & (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ) & (\a[19]  ^ ~\a[20] )) | ((\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ) & (\a[19]  | \a[20] ) & (~\a[19]  | ~\a[20] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[20]  & \b[0]  & (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ));
  assign new_n58_ = (~\b[0]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[1]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[17]  & (~\b[0]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[0]  | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[1]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[2]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & \b[0]  & (~\a[17]  | ~\a[18] ) & (\a[17]  | \a[18] );
  assign new_n59_ = \a[17]  ^ (((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[2]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[3]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )));
  assign new_n60_ = ((~\b[0]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[1]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[17]  & (~\b[0]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[0]  | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[1]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[2]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))) ^ (\b[0]  & (~\a[17]  | ~\a[18] ) & (\a[17]  | \a[18] ));
  assign new_n61_ = \a[14]  ^ (((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n62_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[9]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  ^ \a[14] )) & (~\b[7]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n62_ = (~\b[6]  | ~\b[7] ) & ((\b[6]  & \b[7] ) | (~\b[6]  & ~\b[7] ) | ((~\b[5]  | ~\b[6] ) & ((\b[5]  & \b[6] ) | (~\b[5]  & ~\b[6] ) | ((~\b[4]  | ~\b[5] ) & (((~\b[3]  | ~\b[4] ) & ((\b[3]  & \b[4] ) | (~\b[3]  & ~\b[4] ) | ((~\b[2]  | ~\b[3] ) & ((~\b[2]  & ~\b[3] ) | (\b[2]  & \b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] ))))) | (\b[4]  & \b[5] ) | (~\b[4]  & ~\b[5] ))))));
  assign new_n63_ = ((~\b[0]  | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[1]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[2]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))) ^ (~\a[20]  | ((~\b[0]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[1]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[20]  & (~\b[0]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ))));
  assign new_n64_ = (new_n65_ | ~new_n67_) & ((~new_n65_ & new_n67_) | (new_n65_ & ~new_n67_) | ((~new_n68_ | new_n69_) & (((new_n70_ | ~new_n78_) & (new_n71_ | (~new_n70_ & new_n78_) | (new_n70_ & ~new_n78_))) | (new_n68_ & ~new_n69_) | (~new_n68_ & new_n69_))));
  assign new_n65_ = \a[14]  ^ ((~new_n66_ | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & (~\b[6]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[7]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  ^ \a[14] )) & (~\b[5]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n66_ = (\b[6]  ^ \b[7] ) ^ ((\b[5]  & \b[6] ) | ((~\b[5]  | ~\b[6] ) & (\b[5]  | \b[6] ) & ((\b[4]  & \b[5] ) | (((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))) & (~\b[4]  | ~\b[5] ) & (\b[4]  | \b[5] )))));
  assign new_n67_ = (new_n58_ | (~new_n59_ & new_n60_)) ^ (new_n57_ ^ (~\a[17]  ^ (new_n56_ & (~new_n54_ | ~new_n55_))));
  assign new_n68_ = ~new_n59_ ^ new_n60_;
  assign new_n69_ = \a[14]  ^ ((~new_n50_ | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & (~\b[5]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[6]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  ^ \a[14] )) & (~\b[4]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n70_ = \a[14]  ^ ((~new_n52_ | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & (~\b[4]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[5]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  ^ \a[14] )) & (~\b[3]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n71_ = (~new_n74_ | (\a[14]  ^ (new_n73_ & (~new_n55_ | ~new_n72_)))) & ((~new_n75_ & (new_n76_ | ~new_n77_)) | (new_n74_ & (~\a[14]  ^ (new_n73_ & (~new_n55_ | ~new_n72_)))) | (~new_n74_ & (~\a[14]  | ~new_n73_ | (new_n55_ & new_n72_)) & (\a[14]  | (new_n73_ & (~new_n55_ | ~new_n72_)))));
  assign new_n72_ = (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ) & (\a[13]  | \a[14] ) & (~\a[13]  | ~\a[14] );
  assign new_n73_ = (~\b[3]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[4]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & (~\b[2]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ));
  assign new_n74_ = ((\b[0]  & (\a[15]  | \a[16] ) & (~\a[15]  | ~\a[16] ) & (\a[14]  ^ ~\a[15] )) | (\b[1]  & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ) & (\a[16]  ^ ~\a[17] )) | ((\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ) & (\a[16]  | \a[17] ) & (~\a[16]  | ~\a[17] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[17]  & \b[0]  & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ));
  assign new_n75_ = \b[0]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] ) & (~\b[0]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[1]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[1]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[2]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ));
  assign new_n76_ = \a[14]  ^ (((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[3]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & (~\b[1]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] )));
  assign new_n77_ = (\b[0]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) ^ ((~\b[0]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[1]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[1]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[2]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] )));
  assign new_n78_ = ((~\b[0]  | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[1]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[2]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))) ^ (~\a[17]  | ((~\b[0]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[1]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[17]  & (~\b[0]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ))));
  assign new_n79_ = ~new_n61_ ^ ((~new_n46_ ^ new_n49_) ^ ((~new_n51_ & new_n63_) | (~new_n53_ & (new_n51_ | ~new_n63_) & (~new_n51_ | new_n63_))));
  assign new_n80_ = ~new_n87_ ^ ((~new_n81_ ^ new_n82_) ^ ((new_n46_ & ~new_n49_) | ((~new_n46_ | new_n49_) & (new_n46_ | ~new_n49_) & ((~new_n51_ & new_n63_) | (~new_n53_ & (new_n51_ | ~new_n63_) & (~new_n51_ | new_n63_))))));
  assign new_n81_ = \a[17]  ^ ((~new_n66_ | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )) & (~\b[5]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & (~\b[6]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[7]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  ^ \a[17] )));
  assign new_n82_ = (new_n86_ | (~new_n47_ & new_n48_)) ^ (~new_n85_ ^ (~\a[20]  ^ (new_n84_ & (~new_n83_ | ~new_n55_))));
  assign new_n83_ = (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ) & (\a[19]  | \a[20] ) & (~\a[19]  | ~\a[20] );
  assign new_n84_ = (~\b[2]  | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[3]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[4]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] ));
  assign new_n85_ = (~\b[0]  | ~\a[21]  | (~\a[20]  & \a[21] ) | (\a[20]  & ~\a[21] )) & (~\b[1]  | (~\a[20]  ^ \a[21] ));
  assign new_n86_ = \b[0]  & (\a[20]  ^ \a[21] ) & (~\b[0]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[1]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[20]  & (~\b[0]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[0]  | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[1]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[2]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )));
  assign new_n87_ = \a[14]  ^ (new_n88_ & (~new_n72_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n62_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n88_ = (~\b[9]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[10]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & (~\b[8]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ));
  assign new_n89_ = \a[14]  ^ ((~\b[7]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[8]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  ^ \a[14] )) & (~\b[6]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n62_ & (~\b[7]  ^ \b[8] ))));
  assign new_n90_ = ~new_n91_ & (~new_n79_ | ((new_n89_ | (~new_n53_ & (~new_n51_ | new_n63_) & (new_n51_ | ~new_n63_)) | (new_n53_ & (~new_n51_ ^ ~new_n63_))) & (new_n64_ | (~new_n89_ & (new_n53_ | (new_n51_ & ~new_n63_) | (~new_n51_ & new_n63_)) & (~new_n53_ | (new_n51_ ^ ~new_n63_))) | (new_n89_ & (new_n53_ ^ (new_n51_ ^ ~new_n63_)))))) & (new_n79_ | (~new_n89_ & (new_n53_ | (new_n51_ & ~new_n63_) | (~new_n51_ & new_n63_)) & (~new_n53_ | (new_n51_ ^ ~new_n63_))) | (~new_n64_ & (new_n89_ | (~new_n53_ & (~new_n51_ | new_n63_) & (new_n51_ | ~new_n63_)) | (new_n53_ & (~new_n51_ ^ ~new_n63_))) & (~new_n89_ | (~new_n53_ ^ (new_n51_ ^ ~new_n63_)))));
  assign new_n91_ = \a[11]  ^ (((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~new_n92_ ^ ~\b[11] )) & (~\b[11]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[10]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n92_ = (~\b[10]  | ~\b[11] ) & ((\b[10]  & \b[11] ) | (~\b[10]  & ~\b[11] ) | ((~\b[9]  | ~\b[10] ) & ((\b[9]  & \b[10] ) | (~\b[9]  & ~\b[10] ) | ((~\b[8]  | ~\b[9] ) & ((~\b[8]  & ~\b[9] ) | (\b[8]  & \b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n62_ | (~\b[7]  & ~\b[8] ) | (\b[7]  & \b[8] ))))))));
  assign new_n93_ = ~new_n95_ & (new_n64_ | ~new_n94_) & (~new_n64_ | new_n94_);
  assign new_n94_ = ~new_n89_ ^ (~new_n53_ ^ (~new_n51_ ^ new_n63_));
  assign new_n95_ = \a[11]  ^ ((~new_n96_ | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[10]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[11]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[9]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n96_ = (\b[10]  ^ \b[11] ) ^ ((\b[9]  & \b[10] ) | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((\b[8]  | \b[9] ) & (~\b[8]  | ~\b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (\b[7]  | \b[8] ) & (~\b[7]  | ~\b[8] )))))));
  assign new_n97_ = (~new_n99_ | new_n117_) & ((~new_n100_ & (~new_n116_ | ((new_n119_ | (new_n98_ & ~new_n71_) | (~new_n98_ & new_n71_)) & (new_n102_ | (~new_n119_ & (~new_n98_ | new_n71_) & (new_n98_ | ~new_n71_)) | (new_n119_ & (~new_n98_ ^ ~new_n71_)))))) | (new_n99_ & ~new_n117_) | (~new_n99_ & new_n117_));
  assign new_n98_ = ~new_n70_ ^ new_n78_;
  assign new_n99_ = (~new_n65_ ^ new_n67_) ^ ((new_n68_ & ~new_n69_) | (((~new_n70_ & new_n78_) | (~new_n71_ & (new_n70_ | ~new_n78_) & (~new_n70_ | new_n78_))) & (~new_n68_ | new_n69_) & (new_n68_ | ~new_n69_)));
  assign new_n100_ = ~new_n101_ & ((~new_n68_ & new_n69_) | (new_n68_ & ~new_n69_) | ((new_n70_ | ~new_n78_) & (new_n71_ | (~new_n70_ & new_n78_) | (new_n70_ & ~new_n78_)))) & ((~new_n68_ ^ new_n69_) | (~new_n70_ & new_n78_) | (~new_n71_ & (new_n70_ | ~new_n78_) & (~new_n70_ | new_n78_)));
  assign new_n101_ = \a[11]  ^ (((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n62_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[9]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[7]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n102_ = (new_n103_ | ~new_n104_) & ((~new_n103_ & new_n104_) | (new_n103_ & ~new_n104_) | ((~new_n105_ | new_n106_) & (((new_n107_ | ~new_n115_) & (new_n108_ | (~new_n107_ & new_n115_) | (new_n107_ & ~new_n115_))) | (new_n105_ & ~new_n106_) | (~new_n105_ & new_n106_))));
  assign new_n103_ = \a[11]  ^ ((~new_n66_ | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[6]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[7]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[5]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n104_ = (new_n75_ | (~new_n76_ & new_n77_)) ^ (new_n74_ ^ (~\a[14]  ^ (new_n73_ & (~new_n55_ | ~new_n72_))));
  assign new_n105_ = ~new_n76_ ^ new_n77_;
  assign new_n106_ = \a[11]  ^ ((~new_n50_ | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[5]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[6]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[4]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n107_ = \a[11]  ^ ((~new_n52_ | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[4]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[5]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[3]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n108_ = (~new_n111_ | (\a[11]  ^ (new_n110_ & (~new_n55_ | ~new_n109_)))) & ((~new_n112_ & (new_n113_ | ~new_n114_)) | (new_n111_ & (~\a[11]  ^ (new_n110_ & (~new_n55_ | ~new_n109_)))) | (~new_n111_ & (~\a[11]  | ~new_n110_ | (new_n55_ & new_n109_)) & (\a[11]  | (new_n110_ & (~new_n55_ | ~new_n109_)))));
  assign new_n109_ = (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] );
  assign new_n110_ = (~\b[3]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[4]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[2]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ));
  assign new_n111_ = ((\b[0]  & (\a[12]  | \a[13] ) & (~\a[12]  | ~\a[13] ) & (\a[11]  ^ ~\a[12] )) | (\b[1]  & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ) & (\a[13]  ^ ~\a[14] )) | ((\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ) & (\a[13]  | \a[14] ) & (~\a[13]  | ~\a[14] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[14]  & \b[0]  & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ));
  assign new_n112_ = \b[0]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] ) & (~\b[0]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[1]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[1]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[2]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ));
  assign new_n113_ = \a[11]  ^ (((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[3]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[1]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] )));
  assign new_n114_ = (\b[0]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] )) ^ ((~\b[0]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[1]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[1]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[2]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] )));
  assign new_n115_ = (~\a[14]  | ((~\b[0]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[1]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )))) ^ ((~\b[1]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[2]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] )));
  assign new_n116_ = ~new_n101_ ^ ((~new_n68_ ^ new_n69_) ^ ((~new_n70_ & new_n78_) | (~new_n71_ & (new_n70_ | ~new_n78_) & (~new_n70_ | new_n78_))));
  assign new_n117_ = \a[11]  ^ (new_n118_ & (~new_n109_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n62_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n118_ = (~\b[9]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[10]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[8]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ));
  assign new_n119_ = \a[11]  ^ ((~\b[7]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[8]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[6]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n62_ & (~\b[7]  ^ \b[8] ))));
  assign new_n120_ = ~new_n95_ ^ (~new_n64_ ^ new_n94_);
  assign new_n121_ = ~new_n91_ ^ (new_n79_ ^ ((~new_n89_ & (new_n53_ | (new_n51_ & ~new_n63_) | (~new_n51_ & new_n63_)) & (~new_n53_ | (new_n51_ ^ ~new_n63_))) | (~new_n64_ & (new_n89_ | (~new_n53_ & (~new_n51_ | new_n63_) & (new_n51_ | ~new_n63_)) | (new_n53_ & (~new_n51_ ^ ~new_n63_))) & (~new_n89_ | (~new_n53_ ^ (new_n51_ ^ ~new_n63_))))));
  assign new_n122_ = \a[11]  ^ (~\b[11]  | (((~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (new_n92_ | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ))));
  assign new_n123_ = ~new_n141_ ^ (new_n135_ ^ ((new_n124_ & ~new_n142_) | ((~new_n124_ | new_n142_) & (new_n124_ | ~new_n142_) & (new_n131_ | (~new_n133_ & new_n134_)))));
  assign new_n124_ = new_n129_ ^ (new_n125_ | (~new_n127_ & new_n128_));
  assign new_n125_ = ((\b[2]  & (\a[20]  ^ \a[21] )) | (\b[1]  & \a[21]  & (\a[20]  | ~\a[21] ) & (~\a[20]  | \a[21] ))) & (~\a[20]  ^ (new_n126_ & (~new_n83_ | ~new_n52_)));
  assign new_n126_ = (~\b[3]  | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[4]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[5]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] ));
  assign new_n127_ = (new_n85_ | (\a[20]  ^ (new_n84_ & (~new_n83_ | ~new_n55_)))) & ((~new_n86_ & (new_n47_ | ~new_n48_)) | (~new_n85_ & (~\a[20]  ^ (new_n84_ & (~new_n83_ | ~new_n55_)))) | (new_n85_ & (~\a[20]  | ~new_n84_ | (new_n83_ & new_n55_)) & (\a[20]  | (new_n84_ & (~new_n83_ | ~new_n55_)))));
  assign new_n128_ = ((\b[2]  & (\a[20]  ^ \a[21] )) | (\b[1]  & \a[21]  & (\a[20]  | ~\a[21] ) & (~\a[20]  | \a[21] ))) ^ (~\a[20]  ^ (new_n126_ & (~new_n83_ | ~new_n52_)));
  assign new_n129_ = ((\b[3]  & (\a[20]  ^ \a[21] )) | (\b[2]  & \a[21]  & (\a[20]  | ~\a[21] ) & (~\a[20]  | \a[21] ))) ^ (~\a[20]  ^ (new_n130_ & (~new_n83_ | ~new_n50_)));
  assign new_n130_ = (~\b[4]  | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[5]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[6]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] ));
  assign new_n131_ = ~new_n132_ & (new_n127_ | ~new_n128_) & (~new_n127_ | new_n128_);
  assign new_n132_ = \a[17]  ^ ((~\b[6]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & (~\b[7]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[8]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  ^ \a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n62_ & (~\b[7]  ^ \b[8] ))));
  assign new_n133_ = (new_n81_ | ~new_n82_) & ((~new_n81_ & new_n82_) | (new_n81_ & ~new_n82_) | ((~new_n46_ | new_n49_) & (((new_n51_ | ~new_n63_) & (new_n53_ | (~new_n51_ & new_n63_) | (new_n51_ & ~new_n63_))) | (new_n46_ & ~new_n49_) | (~new_n46_ & new_n49_))));
  assign new_n134_ = ~new_n132_ ^ (~new_n127_ ^ new_n128_);
  assign new_n135_ = ~new_n139_ ^ (new_n137_ ^ (new_n136_ | (new_n129_ & (new_n125_ | (~new_n127_ & new_n128_)))));
  assign new_n136_ = ((\b[3]  & (\a[20]  ^ \a[21] )) | (\b[2]  & \a[21]  & (\a[20]  | ~\a[21] ) & (~\a[20]  | \a[21] ))) & (~\a[20]  ^ (new_n130_ & (~new_n83_ | ~new_n50_)));
  assign new_n137_ = ((\b[4]  & (\a[20]  ^ \a[21] )) | (\b[3]  & \a[21]  & (\a[20]  | ~\a[21] ) & (~\a[20]  | \a[21] ))) ^ (~\a[20]  ^ (new_n138_ & (~new_n83_ | ~new_n66_)));
  assign new_n138_ = (~\b[5]  | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[6]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[7]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] ));
  assign new_n139_ = \a[17]  ^ (new_n140_ & (~new_n54_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n62_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n140_ = (~\b[8]  | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[9]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[10]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] ));
  assign new_n141_ = \a[14]  ^ (~\b[11]  | (((~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & (new_n92_ | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ))));
  assign new_n142_ = \a[17]  ^ ((~\b[7]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & (~\b[8]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[9]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  ^ \a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n62_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))));
  assign new_n143_ = ~new_n144_ & ((new_n124_ & ~new_n142_) | (~new_n124_ & new_n142_) | (~new_n131_ & (new_n133_ | ~new_n134_))) & ((new_n124_ ^ ~new_n142_) | new_n131_ | (~new_n133_ & new_n134_));
  assign new_n144_ = \a[14]  ^ (((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~new_n92_ ^ ~\b[11] )) & (~\b[11]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[10]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n145_ = ~new_n133_ ^ new_n134_;
  assign new_n146_ = (~new_n148_ | new_n87_) & ((~new_n45_ & (~new_n79_ | ((new_n89_ | (new_n147_ & ~new_n53_) | (~new_n147_ & new_n53_)) & (new_n64_ | (~new_n89_ & (~new_n147_ | new_n53_) & (new_n147_ | ~new_n53_)) | (new_n89_ & (~new_n147_ ^ ~new_n53_)))))) | (new_n148_ & ~new_n87_) | (~new_n148_ & new_n87_));
  assign new_n147_ = ~new_n51_ ^ new_n63_;
  assign new_n148_ = (~new_n81_ ^ new_n82_) ^ ((new_n46_ & ~new_n49_) | (((~new_n51_ & new_n63_) | (~new_n53_ & (new_n51_ | ~new_n63_) & (~new_n51_ | new_n63_))) & (~new_n46_ | new_n49_) & (new_n46_ | ~new_n49_)));
  assign new_n149_ = ~new_n144_ ^ ((new_n124_ ^ ~new_n142_) ^ (new_n131_ | (~new_n133_ & new_n134_)));
  assign new_n150_ = \a[14]  ^ ((~new_n96_ | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & (~\b[10]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[11]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  ^ \a[14] )) & (~\b[9]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n151_ = new_n166_ ^ (new_n152_ | (new_n165_ & ((~new_n172_ & new_n173_) | (~new_n163_ & (new_n172_ | ~new_n173_) & (~new_n172_ | new_n173_)))));
  assign new_n152_ = ~new_n153_ & (~new_n159_ | (~new_n154_ & ~new_n162_)) & (new_n159_ | new_n154_ | new_n162_);
  assign new_n153_ = \a[17]  ^ (((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~new_n92_ ^ ~\b[11] )) & (~\b[10]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & (~\b[11]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )));
  assign new_n154_ = new_n156_ & (new_n155_ | (new_n137_ & (new_n136_ | (new_n129_ & (new_n125_ | (~new_n127_ & new_n128_))))));
  assign new_n155_ = ((\b[4]  & (\a[20]  ^ \a[21] )) | (\b[3]  & \a[21]  & (\a[20]  | ~\a[21] ) & (~\a[20]  | \a[21] ))) & (~\a[20]  ^ (new_n138_ & (~new_n83_ | ~new_n66_)));
  assign new_n156_ = ~new_n157_ ^ (~\a[20]  ^ (new_n158_ & (~new_n83_ | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n62_ & (~\b[7]  ^ \b[8] )))));
  assign new_n157_ = (~\b[4]  | ~\a[21]  | (~\a[20]  & \a[21] ) | (\a[20]  & ~\a[21] )) & (~\b[5]  | (~\a[20]  ^ \a[21] ));
  assign new_n158_ = (~\b[6]  | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[7]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[8]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] ));
  assign new_n159_ = ~new_n160_ ^ ~new_n161_;
  assign new_n160_ = \a[20]  ^ ((~\b[7]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  ^ ~\a[19] )) & (~\b[8]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[9]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  ^ \a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n62_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))));
  assign new_n161_ = (~\b[5]  | ~\a[21]  | (~\a[20]  & \a[21] ) | (\a[20]  & ~\a[21] )) & (~\b[6]  | (~\a[20]  ^ \a[21] ));
  assign new_n162_ = ~new_n157_ & (~\a[20]  ^ (new_n158_ & (~new_n83_ | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n62_ & (~\b[7]  ^ \b[8] )))));
  assign new_n163_ = (~new_n164_ | new_n139_) & ((new_n164_ & ~new_n139_) | (~new_n164_ & new_n139_) | ((~new_n124_ | new_n142_) & ((~new_n131_ & (new_n133_ | ~new_n134_)) | (new_n124_ & ~new_n142_) | (~new_n124_ & new_n142_))));
  assign new_n164_ = new_n137_ ^ (new_n136_ | (new_n129_ & (new_n125_ | (~new_n127_ & new_n128_))));
  assign new_n165_ = ~new_n153_ ^ (new_n159_ ^ (new_n154_ | new_n162_));
  assign new_n166_ = ~new_n171_ ^ (new_n167_ ^ ((~new_n160_ & ~new_n161_) | ((~new_n160_ | ~new_n161_) & (new_n160_ | new_n161_) & (new_n154_ | new_n162_))));
  assign new_n167_ = ~new_n170_ ^ (new_n168_ ^ ~\a[20] );
  assign new_n168_ = new_n169_ & (~new_n83_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n62_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))))));
  assign new_n169_ = (~\b[8]  | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[9]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[10]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] ));
  assign new_n170_ = (~\b[6]  | ~\a[21]  | (~\a[20]  & \a[21] ) | (\a[20]  & ~\a[21] )) & (~\b[7]  | (~\a[20]  ^ \a[21] ));
  assign new_n171_ = \a[17]  ^ (~\b[11]  | (((\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & (new_n92_ | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ))));
  assign new_n172_ = \a[17]  ^ ((~new_n96_ | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )) & (~\b[9]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & (~\b[10]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[11]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  ^ \a[17] )));
  assign new_n173_ = new_n156_ ^ (new_n155_ | (new_n137_ & (new_n136_ | (new_n129_ & (new_n125_ | (~new_n127_ & new_n128_))))));
  assign new_n174_ = new_n165_ ^ ((~new_n172_ & new_n173_) | (~new_n163_ & (~new_n172_ | new_n173_) & (new_n172_ | ~new_n173_)));
  assign new_n175_ = ~new_n176_ & (~new_n123_ | (~new_n143_ & (~new_n149_ | ((~new_n145_ | new_n150_) & (new_n146_ | (new_n145_ & ~new_n150_) | (~new_n145_ & new_n150_))))));
  assign new_n176_ = ~new_n141_ & (~new_n135_ | ((~new_n124_ | new_n142_) & ((new_n124_ & ~new_n142_) | (~new_n124_ & new_n142_) | (~new_n131_ & (new_n133_ | ~new_n134_))))) & (new_n135_ | (new_n124_ & ~new_n142_) | ((~new_n124_ | new_n142_) & (new_n124_ | ~new_n142_) & (new_n131_ | (~new_n133_ & new_n134_))));
  assign new_n177_ = ~new_n172_ ^ new_n173_;
  assign new_n178_ = ~new_n179_ ^ (\a[14]  ^ ((new_n190_ ^ \a[17] ) ^ ((\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~new_n189_ & (~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (\a[17]  | (~new_n194_ ^ new_n186_))))));
  assign new_n179_ = (~new_n182_ | ~\a[14] ) & ((new_n182_ & \a[14] ) | (~new_n182_ & ~\a[14] ) | ((~new_n151_ | ~\a[14] ) & ((~new_n151_ & ~\a[14] ) | (new_n151_ & \a[14] ) | ((~new_n174_ | ~\a[14] ) & ((~new_n180_ & (new_n175_ | ~new_n181_)) | (new_n174_ & \a[14] ) | (~new_n174_ & ~\a[14] ))))));
  assign new_n180_ = \a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_);
  assign new_n181_ = \a[14]  ^ (~new_n163_ ^ new_n177_);
  assign new_n182_ = new_n184_ ^ (new_n183_ | (new_n166_ & (new_n152_ | (new_n165_ & ((~new_n172_ & new_n173_) | (~new_n163_ & (new_n172_ | ~new_n173_) & (~new_n172_ | new_n173_)))))));
  assign new_n183_ = ~new_n171_ & (~new_n167_ | ((new_n160_ | new_n161_) & ((new_n160_ & new_n161_) | (~new_n160_ & ~new_n161_) | (~new_n154_ & ~new_n162_)))) & (new_n167_ | (~new_n160_ & ~new_n161_) | ((~new_n160_ | ~new_n161_) & (new_n160_ | new_n161_) & (new_n154_ | new_n162_)));
  assign new_n184_ = \a[17]  ^ (new_n186_ ^ ((~new_n185_ & ~new_n170_) | (((~new_n160_ & ~new_n161_) | ((~new_n160_ | ~new_n161_) & (new_n160_ | new_n161_) & (new_n154_ | new_n162_))) & (~new_n185_ | ~new_n170_) & (new_n185_ | new_n170_))));
  assign new_n185_ = ~new_n168_ ^ ~\a[20] ;
  assign new_n186_ = (new_n187_ ^ ~\a[20] ) ^ ((\b[8]  & (\a[20]  ^ \a[21] )) | (\b[7]  & \a[21]  & (\a[20]  | ~\a[21] ) & (~\a[20]  | \a[21] )));
  assign new_n187_ = new_n188_ & (~new_n83_ | ((~\b[10]  | ~\b[11] ) & (\b[10]  | \b[11] ) & ((\b[9]  & \b[10] ) | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))))) | ((~\b[10]  ^ \b[11] ) & (~\b[9]  | ~\b[10] ) & ((\b[9]  & \b[10] ) | (~\b[9]  & ~\b[10] ) | ((~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n62_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))))))));
  assign new_n188_ = (~\b[9]  | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[10]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[11]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] ));
  assign new_n189_ = ~new_n183_ & (~new_n166_ | (~new_n152_ & (~new_n165_ | ((new_n172_ | ~new_n173_) & (new_n163_ | (~new_n172_ & new_n173_) | (new_n172_ & ~new_n173_))))));
  assign new_n190_ = ~new_n191_ ^ ((new_n193_ ^ ~\a[20] ) ^ ((\b[9]  & (~\a[20]  ^ ~\a[21] )) | (\b[8]  & \a[21]  & (~\a[20]  | \a[21] ) & (\a[20]  | ~\a[21] ))));
  assign new_n191_ = ~new_n192_ & (~new_n186_ | ((new_n185_ | new_n170_) & ((new_n185_ & new_n170_) | (~new_n185_ & ~new_n170_) | ((new_n160_ | new_n161_) & ((new_n160_ & new_n161_) | (~new_n160_ & ~new_n161_) | (~new_n154_ & ~new_n162_))))));
  assign new_n192_ = (new_n187_ ^ ~\a[20] ) & ((\b[8]  & (\a[20]  ^ \a[21] )) | (\b[7]  & \a[21]  & (\a[20]  | ~\a[21] ) & (~\a[20]  | \a[21] )));
  assign new_n193_ = ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~new_n92_ ^ ~\b[11] )) & (~\b[10]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  ^ ~\a[19] )) & (~\b[11]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ));
  assign new_n194_ = (new_n185_ | new_n170_) & (~new_n167_ | ((new_n160_ | new_n161_) & ((new_n160_ & new_n161_) | (~new_n160_ & ~new_n161_) | (~new_n154_ & ~new_n162_))));
  assign new_n195_ = ((\a[11]  & (((~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (new_n175_ | (\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~\a[14]  & (new_n163_ ^ new_n177_)))) | (new_n174_ & \a[14] ) | (~new_n174_ & ~\a[14] )) & ((\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~new_n175_ & (~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (\a[14]  | (~new_n163_ ^ new_n177_))) | (new_n174_ ^ \a[14] ))) | (((\a[11]  & (new_n175_ | (\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~\a[14]  & (new_n163_ ^ new_n177_))) & (~new_n175_ | (\a[14]  ^ (~new_n163_ ^ new_n177_)))) | (~new_n42_ & (~\a[11]  | (~new_n175_ & (~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (\a[14]  | (~new_n163_ ^ new_n177_))) | (new_n175_ & (~\a[14]  ^ (~new_n163_ ^ new_n177_)))) & (\a[11]  | (~new_n175_ ^ (\a[14]  ^ (~new_n163_ ^ new_n177_)))))) & (~\a[11]  | (((\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~new_n175_ & (~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (\a[14]  | (~new_n163_ ^ new_n177_)))) & (~new_n174_ | ~\a[14] ) & (new_n174_ | \a[14] )) | ((~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (new_n175_ | (\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~\a[14]  & (new_n163_ ^ new_n177_))) & (~new_n174_ ^ \a[14] ))) & (\a[11]  | (((\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~new_n175_ & (~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (\a[14]  | (~new_n163_ ^ new_n177_)))) ^ (new_n174_ ^ \a[14] ))))) ^ (\a[11]  ^ ((new_n151_ ^ \a[14] ) ^ ((new_n174_ & \a[14] ) | (((\a[14]  & (new_n163_ | ~new_n177_) & (~new_n163_ | new_n177_)) | (~new_n175_ & (~\a[14]  | (~new_n163_ & new_n177_) | (new_n163_ & ~new_n177_)) & (\a[14]  | (~new_n163_ ^ new_n177_)))) & (~new_n174_ | ~\a[14] ) & (new_n174_ | \a[14] )))));
  assign new_n196_ = new_n198_ ^ ((new_n197_ & \a[11] ) | (~new_n42_ & (new_n197_ | \a[11] ) & (~new_n197_ | ~\a[11] )));
  assign new_n197_ = ~new_n175_ ^ new_n181_;
  assign new_n198_ = \a[11]  ^ ((new_n180_ | (~new_n175_ & new_n181_)) ^ (new_n174_ ^ \a[14] ));
  assign new_n199_ = (~\a[8]  | (~new_n42_ & new_n200_) | (new_n42_ & ~new_n200_)) & (((~new_n201_ | ~\a[8] ) & ((new_n201_ & \a[8] ) | (~new_n201_ & ~\a[8] ) | ((~new_n202_ | ~\a[8] ) & (((~new_n203_ | ~\a[8] ) & (new_n205_ | (new_n203_ & \a[8] ) | (~new_n203_ & ~\a[8] ))) | (new_n202_ & \a[8] ) | (~new_n202_ & ~\a[8] ))))) | (\a[8]  & (new_n42_ | ~new_n200_) & (~new_n42_ | new_n200_)) | (~\a[8]  & (new_n42_ ^ new_n200_)));
  assign new_n200_ = \a[11]  ^ (~new_n175_ ^ new_n181_);
  assign new_n201_ = ((\a[11]  & (~new_n149_ | ((~new_n145_ | new_n150_) & (new_n146_ | (new_n145_ & ~new_n150_) | (~new_n145_ & new_n150_)))) & (new_n149_ | (new_n145_ & ~new_n150_) | (~new_n146_ & (~new_n145_ | new_n150_) & (new_n145_ | ~new_n150_)))) | (((\a[11]  & (new_n146_ | (new_n145_ & ~new_n150_) | (~new_n145_ & new_n150_)) & (~new_n146_ | (new_n145_ ^ ~new_n150_))) | (~new_n43_ & (~\a[11]  | (~new_n146_ & (~new_n145_ | new_n150_) & (new_n145_ | ~new_n150_)) | (new_n146_ & (~new_n145_ ^ ~new_n150_))) & (\a[11]  | (~new_n146_ ^ (new_n145_ ^ ~new_n150_))))) & (~\a[11]  | (new_n149_ & ((new_n145_ & ~new_n150_) | (~new_n146_ & (~new_n145_ | new_n150_) & (new_n145_ | ~new_n150_)))) | (~new_n149_ & (~new_n145_ | new_n150_) & (new_n146_ | (new_n145_ & ~new_n150_) | (~new_n145_ & new_n150_)))) & (\a[11]  | (new_n149_ ^ ((new_n145_ & ~new_n150_) | (~new_n146_ & (~new_n145_ | new_n150_) & (new_n145_ | ~new_n150_))))))) ^ (\a[11]  ^ (new_n123_ ^ (new_n143_ | (new_n149_ & ((new_n145_ & ~new_n150_) | (~new_n146_ & (~new_n145_ | new_n150_) & (new_n145_ | ~new_n150_)))))));
  assign new_n202_ = ((\a[11]  & (new_n146_ | (new_n145_ & ~new_n150_) | (~new_n145_ & new_n150_)) & (~new_n146_ | (new_n145_ ^ ~new_n150_))) | (~new_n43_ & (~\a[11]  | (~new_n146_ & (~new_n145_ | new_n150_) & (new_n145_ | ~new_n150_)) | (new_n146_ & (~new_n145_ ^ ~new_n150_))) & (\a[11]  | (~new_n146_ ^ (new_n145_ ^ ~new_n150_))))) ^ (\a[11]  ^ (new_n149_ ^ ((new_n145_ & ~new_n150_) | (~new_n146_ & (~new_n145_ | new_n150_) & (new_n145_ | ~new_n150_)))));
  assign new_n203_ = ~new_n43_ ^ new_n204_;
  assign new_n204_ = \a[11]  ^ (~new_n146_ ^ (new_n145_ ^ ~new_n150_));
  assign new_n205_ = (~\a[8]  | (new_n206_ & (new_n90_ | (new_n121_ & (new_n93_ | (~new_n97_ & new_n120_))))) | (~new_n206_ & ~new_n90_ & (~new_n121_ | (~new_n93_ & (new_n97_ | ~new_n120_))))) & (((~\a[8]  | (new_n121_ & (new_n93_ | (~new_n97_ & new_n120_))) | (~new_n121_ & ~new_n93_ & (new_n97_ | ~new_n120_))) & (((~\a[8]  | (~new_n97_ & new_n120_) | (new_n97_ & ~new_n120_)) & (new_n207_ | (\a[8]  & (new_n97_ | ~new_n120_) & (~new_n97_ | new_n120_)) | (~\a[8]  & (new_n97_ ^ new_n120_)))) | (\a[8]  & (~new_n121_ | (~new_n93_ & (new_n97_ | ~new_n120_))) & (new_n121_ | new_n93_ | (~new_n97_ & new_n120_))) | (~\a[8]  & (~new_n121_ ^ (new_n93_ | (~new_n97_ & new_n120_)))))) | (\a[8]  & (~new_n206_ | (~new_n90_ & (~new_n121_ | (~new_n93_ & (new_n97_ | ~new_n120_))))) & (new_n206_ | new_n90_ | (new_n121_ & (new_n93_ | (~new_n97_ & new_n120_))))) | (~\a[8]  & (~new_n206_ ^ (new_n90_ | (new_n121_ & (new_n93_ | (~new_n97_ & new_n120_)))))));
  assign new_n206_ = ~new_n44_ ^ new_n122_;
  assign new_n207_ = (~new_n208_ | new_n240_) & ((~new_n210_ & (~new_n239_ | (~new_n212_ & (new_n215_ | ~new_n238_)))) | (new_n208_ & ~new_n240_) | (~new_n208_ & new_n240_));
  assign new_n208_ = new_n209_ ^ (new_n100_ | (new_n116_ & ((~new_n119_ & (new_n71_ | (~new_n70_ & new_n78_) | (new_n70_ & ~new_n78_)) & (~new_n71_ | (~new_n70_ ^ new_n78_))) | (~new_n102_ & (new_n119_ | (~new_n71_ & (new_n70_ | ~new_n78_) & (~new_n70_ | new_n78_)) | (new_n71_ & (new_n70_ ^ new_n78_))) & (~new_n119_ | (~new_n71_ ^ (~new_n70_ ^ new_n78_)))))));
  assign new_n209_ = ~new_n117_ ^ ((~new_n65_ ^ new_n67_) ^ ((new_n68_ & ~new_n69_) | ((~new_n68_ | new_n69_) & (new_n68_ | ~new_n69_) & ((~new_n70_ & new_n78_) | (~new_n71_ & (new_n70_ | ~new_n78_) & (~new_n70_ | new_n78_))))));
  assign new_n210_ = ~new_n211_ & (~new_n116_ | ((new_n119_ | (~new_n71_ & (~new_n70_ | new_n78_) & (new_n70_ | ~new_n78_)) | (new_n71_ & (~new_n70_ ^ ~new_n78_))) & (new_n102_ | (~new_n119_ & (new_n71_ | (new_n70_ & ~new_n78_) | (~new_n70_ & new_n78_)) & (~new_n71_ | (new_n70_ ^ ~new_n78_))) | (new_n119_ & (new_n71_ ^ (new_n70_ ^ ~new_n78_)))))) & (new_n116_ | (~new_n119_ & (new_n71_ | (new_n70_ & ~new_n78_) | (~new_n70_ & new_n78_)) & (~new_n71_ | (new_n70_ ^ ~new_n78_))) | (~new_n102_ & (new_n119_ | (~new_n71_ & (~new_n70_ | new_n78_) & (new_n70_ | ~new_n78_)) | (new_n71_ & (~new_n70_ ^ ~new_n78_))) & (~new_n119_ | (~new_n71_ ^ (new_n70_ ^ ~new_n78_)))));
  assign new_n211_ = \a[8]  ^ (((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~new_n92_ ^ ~\b[11] )) & (~\b[11]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[10]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n212_ = ~new_n214_ & (new_n102_ | ~new_n213_) & (~new_n102_ | new_n213_);
  assign new_n213_ = ~new_n119_ ^ (~new_n71_ ^ (~new_n70_ ^ new_n78_));
  assign new_n214_ = \a[8]  ^ ((~new_n96_ | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[10]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[11]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[9]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n215_ = (~new_n217_ | new_n235_) & ((~new_n218_ & (~new_n234_ | ((new_n237_ | (new_n216_ & ~new_n108_) | (~new_n216_ & new_n108_)) & (new_n220_ | (~new_n237_ & (~new_n216_ | new_n108_) & (new_n216_ | ~new_n108_)) | (new_n237_ & (~new_n216_ ^ ~new_n108_)))))) | (new_n217_ & ~new_n235_) | (~new_n217_ & new_n235_));
  assign new_n216_ = ~new_n107_ ^ new_n115_;
  assign new_n217_ = (~new_n103_ ^ new_n104_) ^ ((new_n105_ & ~new_n106_) | (((~new_n107_ & new_n115_) | (~new_n108_ & (new_n107_ | ~new_n115_) & (~new_n107_ | new_n115_))) & (~new_n105_ | new_n106_) & (new_n105_ | ~new_n106_)));
  assign new_n218_ = ~new_n219_ & ((~new_n105_ & new_n106_) | (new_n105_ & ~new_n106_) | ((new_n107_ | ~new_n115_) & (new_n108_ | (~new_n107_ & new_n115_) | (new_n107_ & ~new_n115_)))) & ((~new_n105_ ^ new_n106_) | (~new_n107_ & new_n115_) | (~new_n108_ & (new_n107_ | ~new_n115_) & (~new_n107_ | new_n115_)));
  assign new_n219_ = \a[8]  ^ (((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n62_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[9]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[7]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n220_ = (~new_n221_ | new_n222_) & ((~new_n221_ & new_n222_) | (new_n221_ & ~new_n222_) | ((~new_n223_ | new_n224_) & (((new_n225_ | ~new_n233_) & (new_n226_ | (~new_n225_ & new_n233_) | (new_n225_ & ~new_n233_))) | (new_n223_ & ~new_n224_) | (~new_n223_ & new_n224_))));
  assign new_n221_ = (new_n112_ | (~new_n113_ & new_n114_)) ^ (new_n111_ ^ (~\a[11]  ^ (new_n110_ & (~new_n55_ | ~new_n109_))));
  assign new_n222_ = \a[8]  ^ ((~new_n66_ | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[6]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[7]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[5]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n223_ = ~new_n113_ ^ new_n114_;
  assign new_n224_ = \a[8]  ^ ((~new_n50_ | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[5]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[6]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[4]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n225_ = \a[8]  ^ ((~new_n52_ | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[4]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[5]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[3]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n226_ = (~new_n229_ | (\a[8]  ^ (new_n228_ & (~new_n55_ | ~new_n227_)))) & ((~new_n230_ & (new_n231_ | ~new_n232_)) | (new_n229_ & (~\a[8]  ^ (new_n228_ & (~new_n55_ | ~new_n227_)))) | (~new_n229_ & (~\a[8]  | ~new_n228_ | (new_n55_ & new_n227_)) & (\a[8]  | (new_n228_ & (~new_n55_ | ~new_n227_)))));
  assign new_n227_ = (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] );
  assign new_n228_ = (~\b[3]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[4]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[2]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ));
  assign new_n229_ = ((\b[0]  & (\a[9]  | \a[10] ) & (~\a[9]  | ~\a[10] ) & (\a[8]  ^ ~\a[9] )) | (\b[1]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  ^ ~\a[11] )) | ((\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[11]  & \b[0]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ));
  assign new_n230_ = \b[0]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] ) & (~\b[0]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[1]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[1]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[2]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ));
  assign new_n231_ = \a[8]  ^ (((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[3]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[1]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )));
  assign new_n232_ = (\b[0]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] )) ^ ((~\b[0]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[1]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[1]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[2]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )));
  assign new_n233_ = (~\a[11]  | ((~\b[0]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[1]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )))) ^ ((~\b[1]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[2]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] )));
  assign new_n234_ = ~new_n219_ ^ ((~new_n105_ ^ new_n106_) ^ ((~new_n107_ & new_n115_) | (~new_n108_ & (new_n107_ | ~new_n115_) & (~new_n107_ | new_n115_))));
  assign new_n235_ = \a[8]  ^ (new_n236_ & (~new_n227_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n62_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n236_ = (~\b[9]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[10]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[8]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ));
  assign new_n237_ = \a[8]  ^ ((~\b[7]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[8]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[6]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n62_ & (~\b[7]  ^ \b[8] ))));
  assign new_n238_ = ~new_n214_ ^ (~new_n102_ ^ new_n213_);
  assign new_n239_ = ~new_n211_ ^ (new_n116_ ^ ((~new_n119_ & (new_n71_ | (new_n70_ & ~new_n78_) | (~new_n70_ & new_n78_)) & (~new_n71_ | (new_n70_ ^ ~new_n78_))) | (~new_n102_ & (new_n119_ | (~new_n71_ & (~new_n70_ | new_n78_) & (new_n70_ | ~new_n78_)) | (new_n71_ & (~new_n70_ ^ ~new_n78_))) & (~new_n119_ | (~new_n71_ ^ (new_n70_ ^ ~new_n78_))))));
  assign new_n240_ = \a[8]  ^ (~\b[11]  | (((~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (new_n92_ | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ))));
  assign new_n241_ = (new_n182_ ^ \a[14] ) ^ ((new_n151_ & \a[14] ) | ((new_n151_ | \a[14] ) & (~new_n151_ | ~\a[14] ) & ((new_n174_ & \a[14] ) | ((new_n180_ | (~new_n175_ & new_n181_)) & (~new_n174_ | ~\a[14] ) & (new_n174_ | \a[14] )))));
  assign new_n242_ = \a[8]  ^ (((~new_n178_ | ~\a[11] ) & (new_n243_ | (new_n178_ & \a[11] ) | (~new_n178_ & ~\a[11] ))) ^ (~new_n246_ ^ \a[11] ));
  assign new_n243_ = (~new_n241_ | ~\a[11] ) & ((new_n241_ & \a[11] ) | (~new_n241_ & ~\a[11] ) | ((~new_n245_ | ~\a[11] ) & ((new_n245_ & \a[11] ) | (~new_n245_ & ~\a[11] ) | ((~\a[11]  | (new_n244_ & (new_n180_ | (~new_n175_ & new_n181_))) | (~new_n244_ & ~new_n180_ & (new_n175_ | ~new_n181_))) & (((~\a[11]  | (~new_n175_ & new_n181_) | (new_n175_ & ~new_n181_)) & (new_n42_ | (\a[11]  & (new_n175_ | ~new_n181_) & (~new_n175_ | new_n181_)) | (~\a[11]  & (new_n175_ ^ new_n181_)))) | (\a[11]  & (~new_n244_ | (~new_n180_ & (new_n175_ | ~new_n181_))) & (new_n244_ | new_n180_ | (~new_n175_ & new_n181_))) | (~\a[11]  & (~new_n244_ ^ (new_n180_ | (~new_n175_ & new_n181_)))))))));
  assign new_n244_ = ~new_n174_ ^ ~\a[14] ;
  assign new_n245_ = (new_n151_ ^ \a[14] ) ^ ((new_n174_ & \a[14] ) | ((new_n180_ | (~new_n175_ & new_n181_)) & (~new_n174_ | ~\a[14] ) & (new_n174_ | \a[14] )));
  assign new_n246_ = ((~\a[14]  | ((~new_n190_ | ~\a[17] ) & (new_n190_ | \a[17] ) & ((\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~new_n189_ & (~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (\a[17]  | (~new_n194_ ^ new_n186_))))) | ((~new_n190_ ^ \a[17] ) & (~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (new_n189_ | (\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~\a[17]  & (new_n194_ ^ new_n186_))))) & (((~\a[14]  | (~new_n189_ & (~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (\a[17]  | (~new_n194_ ^ new_n186_))) | (new_n189_ & (~\a[17]  ^ (~new_n194_ ^ new_n186_)))) & (new_n247_ | (\a[14]  & (new_n189_ | (\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~\a[17]  & (new_n194_ ^ new_n186_))) & (~new_n189_ | (\a[17]  ^ (~new_n194_ ^ new_n186_)))) | (~\a[14]  & (new_n189_ ^ (\a[17]  ^ (~new_n194_ ^ new_n186_)))))) | (\a[14]  & ((new_n190_ & \a[17] ) | (~new_n190_ & ~\a[17] ) | ((~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (new_n189_ | (\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~\a[17]  & (new_n194_ ^ new_n186_))))) & ((new_n190_ ^ \a[17] ) | (\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~new_n189_ & (~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (\a[17]  | (~new_n194_ ^ new_n186_))))) | (~\a[14]  & ((~new_n190_ ^ \a[17] ) ^ ((\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~new_n189_ & (~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (\a[17]  | (~new_n194_ ^ new_n186_)))))))) ^ (~\a[14]  ^ (((~new_n190_ | ~\a[17] ) & ((new_n190_ & \a[17] ) | (~new_n190_ & ~\a[17] ) | ((~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (new_n189_ | (\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~\a[17]  & (new_n194_ ^ new_n186_)))))) ^ (~new_n248_ ^ \a[17] )));
  assign new_n247_ = (~new_n151_ | ~\a[14] ) & ((new_n151_ & \a[14] ) | (~new_n151_ & ~\a[14] ) | ((~new_n174_ | ~\a[14] ) & ((~new_n180_ & (new_n175_ | ~new_n181_)) | (new_n174_ & \a[14] ) | (~new_n174_ & ~\a[14] ))));
  assign new_n248_ = ((new_n249_ ^ ~\a[20] ) ^ ((~\b[10]  | (~\a[20]  ^ \a[21] )) & (~\b[9]  | ~\a[21]  | (~\a[20]  & \a[21] ) | (\a[20]  & ~\a[21] )))) ^ ((((\b[9]  & (\a[20]  ^ \a[21] )) | (\b[8]  & \a[21]  & (\a[20]  | ~\a[21] ) & (~\a[20]  | \a[21] ))) & (new_n193_ ^ ~\a[20] )) | (~new_n191_ & (((~\b[9]  | (~\a[20]  ^ \a[21] )) & (~\b[8]  | ~\a[21]  | (~\a[20]  & \a[21] ) | (\a[20]  & ~\a[21] ))) | (~new_n193_ ^ ~\a[20] )) & ((\b[9]  & (\a[20]  ^ \a[21] )) | (\b[8]  & \a[21]  & (\a[20]  | ~\a[21] ) & (~\a[20]  | \a[21] )) | (~new_n193_ & ~\a[20] ) | (new_n193_ & \a[20] ))));
  assign new_n249_ = \b[11]  & (((~\a[19]  | ~\a[20] ) & (\a[19]  | \a[20] ) & (\a[17]  ^ ~\a[18] ) & (\a[18]  ^ ~\a[19] )) | (~new_n92_ & (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ) & (~\a[19]  | ~\a[20] ) & (\a[19]  | \a[20] )));
  assign new_n250_ = ((\a[8]  & (new_n41_ | (new_n241_ & \a[11] ) | (~new_n241_ & ~\a[11] )) & (~new_n41_ | (new_n241_ ^ \a[11] ))) | (((new_n195_ & \a[8] ) | ((~new_n195_ | ~\a[8] ) & (new_n195_ | \a[8] ) & ((new_n196_ & \a[8] ) | (~new_n199_ & (~new_n196_ | ~\a[8] ) & (new_n196_ | \a[8] ))))) & (~\a[8]  | (~new_n41_ & (~new_n241_ | ~\a[11] ) & (new_n241_ | \a[11] )) | (new_n41_ & (~new_n241_ ^ \a[11] ))) & (\a[8]  | (~new_n41_ ^ (new_n241_ ^ \a[11] ))))) ^ (\a[8]  ^ ((new_n178_ ^ \a[11] ) ^ ((new_n241_ & \a[11] ) | (~new_n41_ & (~new_n241_ | ~\a[11] ) & (new_n241_ | \a[11] )))));
  assign new_n251_ = ((new_n195_ & \a[8] ) | ((~new_n195_ | ~\a[8] ) & (new_n195_ | \a[8] ) & ((new_n196_ & \a[8] ) | (~new_n199_ & (~new_n196_ | ~\a[8] ) & (new_n196_ | \a[8] ))))) ^ (~new_n252_ ^ ~\a[8] );
  assign new_n252_ = (new_n241_ ^ \a[11] ) ^ ((new_n245_ & \a[11] ) | ((~new_n245_ | ~\a[11] ) & (new_n245_ | \a[11] ) & ((\a[11]  & (~new_n244_ | (~new_n180_ & (new_n175_ | ~new_n181_))) & (new_n244_ | new_n180_ | (~new_n175_ & new_n181_))) | (((\a[11]  & (new_n175_ | ~new_n181_) & (~new_n175_ | new_n181_)) | (~new_n42_ & (~\a[11]  | (~new_n175_ & new_n181_) | (new_n175_ & ~new_n181_)) & (\a[11]  | (~new_n175_ ^ new_n181_)))) & (~\a[11]  | (new_n244_ & (new_n180_ | (~new_n175_ & new_n181_))) | (~new_n244_ & ~new_n180_ & (new_n175_ | ~new_n181_))) & (\a[11]  | (new_n244_ ^ (new_n180_ | (~new_n175_ & new_n181_))))))));
  assign new_n253_ = (~new_n195_ ^ ~\a[8] ) ^ ((new_n196_ & \a[8] ) | (~new_n199_ & (new_n196_ | \a[8] ) & (~new_n196_ | ~\a[8] )));
  assign new_n254_ = (~\a[5]  | (~new_n255_ & new_n199_) | (new_n255_ & ~new_n199_)) & (((~new_n256_ | ~\a[5] ) & ((new_n256_ & \a[5] ) | (~new_n256_ & ~\a[5] ) | ((~new_n257_ | ~\a[5] ) & (((~new_n258_ | ~\a[5] ) & (new_n259_ | (new_n258_ & \a[5] ) | (~new_n258_ & ~\a[5] ))) | (new_n257_ & \a[5] ) | (~new_n257_ & ~\a[5] ))))) | (\a[5]  & (new_n255_ | ~new_n199_) & (~new_n255_ | new_n199_)) | (~\a[5]  & (new_n255_ ^ new_n199_)));
  assign new_n255_ = \a[8]  ^ (new_n198_ ^ ((new_n197_ & \a[11] ) | (~new_n42_ & (new_n197_ | \a[11] ) & (~new_n197_ | ~\a[11] ))));
  assign new_n256_ = ((new_n201_ & \a[8] ) | ((~new_n201_ | ~\a[8] ) & (new_n201_ | \a[8] ) & ((new_n202_ & \a[8] ) | (((new_n203_ & \a[8] ) | (~new_n205_ & (~new_n203_ | ~\a[8] ) & (new_n203_ | \a[8] ))) & (~new_n202_ | ~\a[8] ) & (new_n202_ | \a[8] ))))) ^ (\a[8]  ^ (~new_n42_ ^ new_n200_));
  assign new_n257_ = ((new_n202_ & \a[8] ) | ((~new_n202_ | ~\a[8] ) & (new_n202_ | \a[8] ) & ((new_n203_ & \a[8] ) | (~new_n205_ & (~new_n203_ | ~\a[8] ) & (new_n203_ | \a[8] ))))) ^ (~new_n201_ ^ ~\a[8] );
  assign new_n258_ = (~new_n202_ ^ ~\a[8] ) ^ ((new_n203_ & \a[8] ) | (~new_n205_ & (new_n203_ | \a[8] ) & (~new_n203_ | ~\a[8] )));
  assign new_n259_ = (~\a[5]  | (~new_n205_ & new_n260_) | (new_n205_ & ~new_n260_)) & (((~new_n261_ | ~\a[5] ) & ((new_n261_ & \a[5] ) | (~new_n261_ & ~\a[5] ) | ((~new_n262_ | ~\a[5] ) & (((~new_n263_ | ~\a[5] ) & (new_n265_ | (new_n263_ & \a[5] ) | (~new_n263_ & ~\a[5] ))) | (new_n262_ & \a[5] ) | (~new_n262_ & ~\a[5] ))))) | (\a[5]  & (new_n205_ | ~new_n260_) & (~new_n205_ | new_n260_)) | (~\a[5]  & (new_n205_ ^ new_n260_)));
  assign new_n260_ = \a[8]  ^ (~new_n43_ ^ new_n204_);
  assign new_n261_ = ((\a[8]  & (~new_n121_ | (~new_n93_ & (new_n97_ | ~new_n120_))) & (new_n121_ | new_n93_ | (~new_n97_ & new_n120_))) | (((\a[8]  & (new_n97_ | ~new_n120_) & (~new_n97_ | new_n120_)) | (~new_n207_ & (~\a[8]  | (~new_n97_ & new_n120_) | (new_n97_ & ~new_n120_)) & (\a[8]  | (~new_n97_ ^ new_n120_)))) & (~\a[8]  | (new_n121_ & (new_n93_ | (~new_n97_ & new_n120_))) | (~new_n121_ & ~new_n93_ & (new_n97_ | ~new_n120_))) & (\a[8]  | (new_n121_ ^ (new_n93_ | (~new_n97_ & new_n120_)))))) ^ (\a[8]  ^ (new_n206_ ^ (new_n90_ | (new_n121_ & (new_n93_ | (~new_n97_ & new_n120_))))));
  assign new_n262_ = ((\a[8]  & (~new_n97_ | new_n120_) & (new_n97_ | ~new_n120_)) | (~new_n207_ & (~\a[8]  | (new_n97_ & ~new_n120_) | (~new_n97_ & new_n120_)) & (\a[8]  | (new_n97_ ^ ~new_n120_)))) ^ (\a[8]  ^ (new_n121_ ^ (new_n93_ | (~new_n97_ & new_n120_))));
  assign new_n263_ = ~new_n207_ ^ new_n264_;
  assign new_n264_ = \a[8]  ^ (~new_n97_ ^ new_n120_);
  assign new_n265_ = (~\a[5]  | (new_n266_ & (new_n210_ | (new_n239_ & (new_n212_ | (~new_n215_ & new_n238_))))) | (~new_n266_ & ~new_n210_ & (~new_n239_ | (~new_n212_ & (new_n215_ | ~new_n238_))))) & (((~\a[5]  | (new_n239_ & (new_n212_ | (~new_n215_ & new_n238_))) | (~new_n239_ & ~new_n212_ & (new_n215_ | ~new_n238_))) & (((~\a[5]  | (~new_n215_ & new_n238_) | (new_n215_ & ~new_n238_)) & (new_n267_ | (\a[5]  & (new_n215_ | ~new_n238_) & (~new_n215_ | new_n238_)) | (~\a[5]  & (new_n215_ ^ new_n238_)))) | (\a[5]  & (~new_n239_ | (~new_n212_ & (new_n215_ | ~new_n238_))) & (new_n239_ | new_n212_ | (~new_n215_ & new_n238_))) | (~\a[5]  & (~new_n239_ ^ (new_n212_ | (~new_n215_ & new_n238_)))))) | (\a[5]  & (~new_n266_ | (~new_n210_ & (~new_n239_ | (~new_n212_ & (new_n215_ | ~new_n238_))))) & (new_n266_ | new_n210_ | (new_n239_ & (new_n212_ | (~new_n215_ & new_n238_))))) | (~\a[5]  & (~new_n266_ ^ (new_n210_ | (new_n239_ & (new_n212_ | (~new_n215_ & new_n238_)))))));
  assign new_n266_ = ~new_n208_ ^ new_n240_;
  assign new_n267_ = (~new_n268_ | new_n301_) & ((~new_n270_ & (~new_n300_ | (~new_n272_ & (new_n275_ | ~new_n299_)))) | (new_n268_ & ~new_n301_) | (~new_n268_ & new_n301_));
  assign new_n268_ = new_n269_ ^ (new_n218_ | (new_n234_ & ((~new_n237_ & (new_n108_ | (~new_n107_ & new_n115_) | (new_n107_ & ~new_n115_)) & (~new_n108_ | (~new_n107_ ^ new_n115_))) | (~new_n220_ & (new_n237_ | (~new_n108_ & (new_n107_ | ~new_n115_) & (~new_n107_ | new_n115_)) | (new_n108_ & (new_n107_ ^ new_n115_))) & (~new_n237_ | (~new_n108_ ^ (~new_n107_ ^ new_n115_)))))));
  assign new_n269_ = ~new_n235_ ^ ((~new_n103_ ^ new_n104_) ^ ((new_n105_ & ~new_n106_) | ((~new_n105_ | new_n106_) & (new_n105_ | ~new_n106_) & ((~new_n107_ & new_n115_) | (~new_n108_ & (new_n107_ | ~new_n115_) & (~new_n107_ | new_n115_))))));
  assign new_n270_ = ~new_n271_ & (~new_n234_ | ((new_n237_ | (~new_n108_ & (~new_n107_ | new_n115_) & (new_n107_ | ~new_n115_)) | (new_n108_ & (~new_n107_ ^ ~new_n115_))) & (new_n220_ | (~new_n237_ & (new_n108_ | (new_n107_ & ~new_n115_) | (~new_n107_ & new_n115_)) & (~new_n108_ | (new_n107_ ^ ~new_n115_))) | (new_n237_ & (new_n108_ ^ (new_n107_ ^ ~new_n115_)))))) & (new_n234_ | (~new_n237_ & (new_n108_ | (new_n107_ & ~new_n115_) | (~new_n107_ & new_n115_)) & (~new_n108_ | (new_n107_ ^ ~new_n115_))) | (~new_n220_ & (new_n237_ | (~new_n108_ & (~new_n107_ | new_n115_) & (new_n107_ | ~new_n115_)) | (new_n108_ & (~new_n107_ ^ ~new_n115_))) & (~new_n237_ | (~new_n108_ ^ (new_n107_ ^ ~new_n115_)))));
  assign new_n271_ = \a[5]  ^ (((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~new_n92_ ^ ~\b[11] )) & (~\b[11]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[10]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n272_ = ~new_n274_ & (new_n220_ | ~new_n273_) & (~new_n220_ | new_n273_);
  assign new_n273_ = ~new_n237_ ^ (~new_n108_ ^ (~new_n107_ ^ new_n115_));
  assign new_n274_ = \a[5]  ^ ((~new_n96_ | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[10]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[11]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[9]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n275_ = (~new_n277_ | new_n296_) & ((new_n277_ & ~new_n296_) | (~new_n277_ & new_n296_) | (~new_n278_ & (~new_n280_ | ((new_n298_ | (new_n276_ & ~new_n226_) | (~new_n276_ & new_n226_)) & (new_n281_ | (~new_n298_ & (~new_n276_ | new_n226_) & (new_n276_ | ~new_n226_)) | (new_n298_ & (~new_n276_ ^ ~new_n226_)))))));
  assign new_n276_ = ~new_n225_ ^ new_n233_;
  assign new_n277_ = (~new_n221_ ^ new_n222_) ^ ((new_n223_ & ~new_n224_) | (((~new_n225_ & new_n233_) | (~new_n226_ & (new_n225_ | ~new_n233_) & (~new_n225_ | new_n233_))) & (~new_n223_ | new_n224_) & (new_n223_ | ~new_n224_)));
  assign new_n278_ = ~new_n279_ & ((~new_n223_ & new_n224_) | (new_n223_ & ~new_n224_) | ((new_n225_ | ~new_n233_) & (new_n226_ | (~new_n225_ & new_n233_) | (new_n225_ & ~new_n233_)))) & ((~new_n223_ ^ new_n224_) | (~new_n225_ & new_n233_) | (~new_n226_ & (new_n225_ | ~new_n233_) & (~new_n225_ | new_n233_)));
  assign new_n279_ = \a[5]  ^ (((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n62_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[9]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[7]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n280_ = ~new_n279_ ^ ((~new_n223_ ^ new_n224_) ^ ((~new_n225_ & new_n233_) | (~new_n226_ & (new_n225_ | ~new_n233_) & (~new_n225_ | new_n233_))));
  assign new_n281_ = (~new_n282_ | new_n283_) & ((~new_n282_ & new_n283_) | (new_n282_ & ~new_n283_) | ((~new_n284_ | new_n285_) & (((new_n286_ | ~new_n295_) & (new_n289_ | (~new_n286_ & new_n295_) | (new_n286_ & ~new_n295_))) | (new_n284_ & ~new_n285_) | (~new_n284_ & new_n285_))));
  assign new_n282_ = (new_n230_ | (~new_n231_ & new_n232_)) ^ (new_n229_ ^ (~\a[8]  ^ (new_n228_ & (~new_n55_ | ~new_n227_))));
  assign new_n283_ = \a[5]  ^ ((~new_n66_ | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[6]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[7]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[5]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n284_ = ~new_n231_ ^ new_n232_;
  assign new_n285_ = \a[5]  ^ ((~new_n50_ | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[5]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[6]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[4]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n286_ = \a[5]  ^ (new_n288_ & (~new_n52_ | ~new_n287_));
  assign new_n287_ = (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (\a[4]  | \a[5] ) & (~\a[4]  | ~\a[5] );
  assign new_n288_ = (~\b[4]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[5]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[3]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n289_ = (~new_n291_ | (\a[5]  ^ (new_n290_ & (~new_n55_ | ~new_n287_)))) & ((~new_n292_ & (new_n293_ | ~new_n294_)) | (new_n291_ & (~\a[5]  ^ (new_n290_ & (~new_n55_ | ~new_n287_)))) | (~new_n291_ & (~\a[5]  | ~new_n290_ | (new_n55_ & new_n287_)) & (\a[5]  | (new_n290_ & (~new_n55_ | ~new_n287_)))));
  assign new_n290_ = (~\b[3]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[4]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[2]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n291_ = ((\b[0]  & (\a[6]  | \a[7] ) & (~\a[6]  | ~\a[7] ) & (\a[5]  ^ ~\a[6] )) | (\b[1]  & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (\a[7]  ^ ~\a[8] )) | ((\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[8]  & \b[0]  & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ));
  assign new_n292_ = \b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (~\b[0]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[1]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[1]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[2]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n293_ = \a[5]  ^ (((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[3]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[1]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )));
  assign new_n294_ = (\b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] )) ^ ((~\b[0]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[1]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[1]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[2]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )));
  assign new_n295_ = (~\a[8]  | ((~\b[0]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[1]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )))) ^ ((~\b[1]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[2]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )));
  assign new_n296_ = \a[5]  ^ (new_n297_ & (~new_n287_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n62_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n297_ = (~\b[9]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[10]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[8]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n298_ = \a[5]  ^ ((~\b[7]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[8]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[6]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n62_ & (~\b[7]  ^ \b[8] ))));
  assign new_n299_ = ~new_n274_ ^ (~new_n220_ ^ new_n273_);
  assign new_n300_ = ~new_n271_ ^ (new_n234_ ^ ((~new_n237_ & (new_n108_ | (new_n107_ & ~new_n115_) | (~new_n107_ & new_n115_)) & (~new_n108_ | (new_n107_ ^ ~new_n115_))) | (~new_n220_ & (new_n237_ | (~new_n108_ & (~new_n107_ | new_n115_) & (new_n107_ | ~new_n115_)) | (new_n108_ & (~new_n107_ ^ ~new_n115_))) & (~new_n237_ | (~new_n108_ ^ (new_n107_ ^ ~new_n115_))))));
  assign new_n301_ = \a[5]  ^ (~\b[11]  | (((~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (new_n92_ | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ))));
  assign new_n302_ = (~new_n304_ ^ \a[8] ) ^ ((new_n40_ | ~new_n242_) & (~new_n303_ | ~\a[8] ));
  assign new_n303_ = (new_n246_ ^ ~\a[11] ) ^ ((~new_n178_ | ~\a[11] ) & (new_n243_ | (~new_n178_ & ~\a[11] ) | (new_n178_ & \a[11] )));
  assign new_n304_ = ((new_n246_ & \a[11] ) | (((new_n178_ & \a[11] ) | (~new_n243_ & (~new_n178_ | ~\a[11] ) & (new_n178_ | \a[11] ))) & (~new_n246_ | ~\a[11] ) & (new_n246_ | \a[11] ))) ^ (~\a[11]  ^ (new_n305_ ^ new_n306_));
  assign new_n305_ = (~\a[14]  | ((~new_n190_ | ~\a[17] ) & ((new_n190_ & \a[17] ) | (~new_n190_ & ~\a[17] ) | ((~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (new_n189_ | (\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~\a[17]  & (new_n194_ ^ new_n186_))))) & (~new_n248_ ^ \a[17] )) | (((new_n190_ & \a[17] ) | ((~new_n190_ | ~\a[17] ) & (new_n190_ | \a[17] ) & ((\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~new_n189_ & (~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (\a[17]  | (~new_n194_ ^ new_n186_)))))) & (~new_n248_ | ~\a[17] ) & (new_n248_ | \a[17] ))) & (((~\a[14]  | ((~new_n190_ | ~\a[17] ) & (new_n190_ | \a[17] ) & ((\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~new_n189_ & (~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (\a[17]  | (~new_n194_ ^ new_n186_))))) | ((~new_n190_ ^ \a[17] ) & (~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (new_n189_ | (\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~\a[17]  & (new_n194_ ^ new_n186_))))) & (((~\a[14]  | (~new_n189_ & (~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (\a[17]  | (~new_n194_ ^ new_n186_))) | (new_n189_ & (~\a[17]  ^ (~new_n194_ ^ new_n186_)))) & (new_n247_ | (\a[14]  & (new_n189_ | (\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~\a[17]  & (new_n194_ ^ new_n186_))) & (~new_n189_ | (\a[17]  ^ (~new_n194_ ^ new_n186_)))) | (~\a[14]  & (new_n189_ ^ (\a[17]  ^ (~new_n194_ ^ new_n186_)))))) | (\a[14]  & ((new_n190_ & \a[17] ) | (~new_n190_ & ~\a[17] ) | ((~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (new_n189_ | (\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~\a[17]  & (new_n194_ ^ new_n186_))))) & ((new_n190_ ^ \a[17] ) | (\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~new_n189_ & (~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (\a[17]  | (~new_n194_ ^ new_n186_))))) | (~\a[14]  & ((~new_n190_ ^ \a[17] ) ^ ((\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~new_n189_ & (~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (\a[17]  | (~new_n194_ ^ new_n186_)))))))) | (\a[14]  & ((new_n190_ & \a[17] ) | ((~new_n190_ | ~\a[17] ) & (new_n190_ | \a[17] ) & ((\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~new_n189_ & (~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (\a[17]  | (~new_n194_ ^ new_n186_))))) | (new_n248_ ^ \a[17] )) & (((~new_n190_ | ~\a[17] ) & ((new_n190_ & \a[17] ) | (~new_n190_ & ~\a[17] ) | ((~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (new_n189_ | (\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~\a[17]  & (new_n194_ ^ new_n186_)))))) | (new_n248_ & \a[17] ) | (~new_n248_ & ~\a[17] ))) | (~\a[14]  & (((new_n190_ & \a[17] ) | ((~new_n190_ | ~\a[17] ) & (new_n190_ | \a[17] ) & ((\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~new_n189_ & (~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (\a[17]  | (~new_n194_ ^ new_n186_)))))) ^ (~new_n248_ ^ \a[17] ))));
  assign new_n306_ = \a[14]  ^ ((~new_n307_ ^ \a[17] ) ^ ((~new_n248_ | ~\a[17] ) & (((~new_n190_ | ~\a[17] ) & ((new_n190_ & \a[17] ) | (~new_n190_ & ~\a[17] ) | ((~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (new_n189_ | (\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~\a[17]  & (new_n194_ ^ new_n186_)))))) | (new_n248_ & \a[17] ) | (~new_n248_ & ~\a[17] ))));
  assign new_n307_ = ~new_n308_ ^ (\a[20]  ? ((~\a[21]  | ~\b[10] ) & (~\b[11]  | (~\a[20]  ^ \a[21] ))) : (\a[21]  & \b[11] ));
  assign new_n308_ = ((new_n249_ ^ ~\a[20] ) | ((~\b[10]  | (~\a[20]  ^ \a[21] )) & (~\b[9]  | ~\a[21]  | (~\a[20]  & \a[21] ) | (\a[20]  & ~\a[21] )))) & (((~new_n249_ | \a[20] ) & (new_n249_ | ~\a[20] ) & (~\b[10]  | (~\a[20]  ^ \a[21] )) & (~\b[9]  | ~\a[21]  | (~\a[20]  & \a[21] ) | (\a[20]  & ~\a[21] ))) | ((~new_n249_ ^ ~\a[20] ) & ((\b[10]  & (\a[20]  ^ \a[21] )) | (\b[9]  & \a[21]  & (\a[20]  | ~\a[21] ) & (~\a[20]  | \a[21] )))) | ((((~\b[9]  | (~\a[20]  ^ \a[21] )) & (~\b[8]  | ~\a[21]  | (~\a[20]  & \a[21] ) | (\a[20]  & ~\a[21] ))) | (~new_n193_ ^ ~\a[20] )) & (new_n191_ | (((\b[9]  & (\a[20]  ^ \a[21] )) | (\b[8]  & \a[21]  & (\a[20]  | ~\a[21] ) & (~\a[20]  | \a[21] ))) & (new_n193_ ^ ~\a[20] )) | ((~\b[9]  | (~\a[20]  ^ \a[21] )) & (~\b[8]  | ~\a[21]  | (~\a[20]  & \a[21] ) | (\a[20]  & ~\a[21] )) & (new_n193_ | \a[20] ) & (~new_n193_ | ~\a[20] )))));
  assign new_n309_ = (~\a[2]  | (new_n310_ & ~new_n254_) | (~new_n310_ & new_n254_)) & (((~new_n355_ | ~\a[2] ) & (((~new_n356_ | ~\a[2] ) & (new_n311_ | (new_n356_ & \a[2] ) | (~new_n356_ & ~\a[2] ))) | (new_n355_ & \a[2] ) | (~new_n355_ & ~\a[2] ))) | (\a[2]  & (~new_n310_ | new_n254_) & (new_n310_ | ~new_n254_)) | (~\a[2]  & (~new_n310_ ^ ~new_n254_)));
  assign new_n310_ = ~new_n253_ ^ ~\a[5] ;
  assign new_n311_ = (~\a[2]  | ((~new_n257_ | ~\a[5] ) & (new_n257_ | \a[5] ) & ((new_n258_ & \a[5] ) | ((~new_n258_ | ~\a[5] ) & (new_n258_ | \a[5] ) & ((new_n352_ & \a[5] ) | (~new_n353_ & (~new_n352_ | ~\a[5] ) & (new_n352_ | \a[5] )))))) | ((~new_n257_ ^ \a[5] ) & (~new_n258_ | ~\a[5] ) & ((new_n258_ & \a[5] ) | (~new_n258_ & ~\a[5] ) | ((~new_n352_ | ~\a[5] ) & (new_n353_ | (new_n352_ & \a[5] ) | (~new_n352_ & ~\a[5] )))))) & (((~\a[2]  | ((~new_n258_ | ~\a[5] ) & (new_n258_ | \a[5] ) & ((new_n352_ & \a[5] ) | (~new_n353_ & (~new_n352_ | ~\a[5] ) & (new_n352_ | \a[5] )))) | ((~new_n258_ ^ \a[5] ) & (~new_n352_ | ~\a[5] ) & (new_n353_ | (new_n352_ & \a[5] ) | (~new_n352_ & ~\a[5] )))) & (((~\a[2]  | (~new_n353_ & (~new_n352_ | ~\a[5] ) & (new_n352_ | \a[5] )) | (new_n353_ & (~new_n352_ ^ \a[5] ))) & (((~new_n354_ | ~\a[2] ) & (new_n312_ | (new_n354_ & \a[2] ) | (~new_n354_ & ~\a[2] ))) | (\a[2]  & (new_n353_ | (new_n352_ & \a[5] ) | (~new_n352_ & ~\a[5] )) & (~new_n353_ | (new_n352_ ^ \a[5] ))) | (~\a[2]  & (new_n353_ ^ (new_n352_ ^ \a[5] ))))) | (\a[2]  & ((new_n258_ & \a[5] ) | (~new_n258_ & ~\a[5] ) | ((~new_n352_ | ~\a[5] ) & (new_n353_ | (new_n352_ & \a[5] ) | (~new_n352_ & ~\a[5] )))) & ((new_n258_ ^ \a[5] ) | (new_n352_ & \a[5] ) | (~new_n353_ & (~new_n352_ | ~\a[5] ) & (new_n352_ | \a[5] )))) | (~\a[2]  & ((~new_n258_ ^ \a[5] ) ^ ((new_n352_ & \a[5] ) | (~new_n353_ & (~new_n352_ | ~\a[5] ) & (new_n352_ | \a[5] ))))))) | (\a[2]  & ((new_n257_ & \a[5] ) | (~new_n257_ & ~\a[5] ) | ((~new_n258_ | ~\a[5] ) & ((new_n258_ & \a[5] ) | (~new_n258_ & ~\a[5] ) | ((~new_n352_ | ~\a[5] ) & (new_n353_ | (new_n352_ & \a[5] ) | (~new_n352_ & ~\a[5] )))))) & ((new_n257_ ^ \a[5] ) | (new_n258_ & \a[5] ) | ((~new_n258_ | ~\a[5] ) & (new_n258_ | \a[5] ) & ((new_n352_ & \a[5] ) | (~new_n353_ & (~new_n352_ | ~\a[5] ) & (new_n352_ | \a[5] )))))) | (~\a[2]  & ((~new_n257_ ^ \a[5] ) ^ ((new_n258_ & \a[5] ) | ((~new_n258_ | ~\a[5] ) & (new_n258_ | \a[5] ) & ((new_n352_ & \a[5] ) | (~new_n353_ & (~new_n352_ | ~\a[5] ) & (new_n352_ | \a[5] ))))))));
  assign new_n312_ = (~new_n314_ | ~\a[2] ) & ((new_n314_ & \a[2] ) | (~new_n314_ & ~\a[2] ) | ((~\a[2]  | (~new_n313_ & new_n265_) | (new_n313_ & ~new_n265_)) & (((~new_n350_ | ~\a[2] ) & ((new_n350_ & \a[2] ) | (~new_n350_ & ~\a[2] ) | ((~new_n351_ | ~\a[2] ) & (new_n315_ | (new_n351_ & \a[2] ) | (~new_n351_ & ~\a[2] ))))) | (\a[2]  & (new_n313_ | ~new_n265_) & (~new_n313_ | new_n265_)) | (~\a[2]  & (new_n313_ ^ new_n265_)))));
  assign new_n313_ = ~new_n263_ ^ ~\a[5] ;
  assign new_n314_ = (~new_n262_ ^ ~\a[5] ) ^ ((new_n263_ & \a[5] ) | (~new_n265_ & (new_n263_ | \a[5] ) & (~new_n263_ | ~\a[5] )));
  assign new_n315_ = (~new_n316_ | ~\a[2] ) & ((~new_n316_ & ~\a[2] ) | (new_n316_ & \a[2] ) | ((~new_n348_ | ~\a[2] ) & ((new_n348_ & \a[2] ) | (~new_n348_ & ~\a[2] ) | ((~new_n349_ | ~\a[2] ) & (new_n318_ | (new_n349_ & \a[2] ) | (~new_n349_ & ~\a[2] ))))));
  assign new_n316_ = ~new_n267_ ^ new_n317_;
  assign new_n317_ = \a[5]  ^ (~new_n215_ ^ new_n238_);
  assign new_n318_ = (~\a[2]  | (new_n275_ & ~new_n299_) | (~new_n275_ & new_n299_)) & (((~new_n319_ | new_n347_) & ((new_n319_ & ~new_n347_) | (~new_n319_ & new_n347_) | (~new_n344_ & (new_n321_ | ~new_n346_)))) | (\a[2]  & (~new_n275_ | new_n299_) & (new_n275_ | ~new_n299_)) | (~\a[2]  & (~new_n275_ ^ ~new_n299_)));
  assign new_n319_ = new_n320_ ^ (new_n278_ | (new_n280_ & ((~new_n298_ & (new_n276_ | ~new_n226_) & (~new_n276_ | new_n226_)) | (~new_n281_ & (new_n298_ | (~new_n276_ & new_n226_) | (new_n276_ & ~new_n226_)) & (~new_n298_ | (~new_n276_ ^ new_n226_))))));
  assign new_n320_ = ~new_n277_ ^ new_n296_;
  assign new_n321_ = (new_n338_ | (new_n322_ & ~new_n281_) | (~new_n322_ & new_n281_)) & ((~new_n338_ & (~new_n322_ | new_n281_) & (new_n322_ | ~new_n281_)) | (new_n338_ & (~new_n322_ ^ ~new_n281_)) | ((~new_n339_ | new_n343_) & ((~new_n339_ & new_n343_) | (new_n339_ & ~new_n343_) | (~new_n340_ & (new_n323_ | ~new_n342_)))));
  assign new_n322_ = ~new_n298_ ^ (~new_n276_ ^ new_n226_);
  assign new_n323_ = (new_n332_ | (new_n324_ & ~new_n289_) | (~new_n324_ & new_n289_)) & ((~new_n332_ & (~new_n324_ | new_n289_) & (new_n324_ | ~new_n289_)) | (new_n332_ & (~new_n324_ ^ ~new_n289_)) | ((new_n333_ | ~new_n334_) & ((~new_n333_ & new_n334_) | (new_n333_ & ~new_n334_) | ((new_n335_ | ~new_n337_) & (new_n325_ | (~new_n335_ & new_n337_) | (new_n335_ & ~new_n337_))))));
  assign new_n324_ = ~new_n286_ ^ new_n295_;
  assign new_n325_ = (~new_n329_ | (\a[2]  ^ (new_n328_ & (~new_n52_ | ~new_n327_)))) & (((new_n326_ | ~new_n330_) & (~new_n331_ | (new_n326_ & ~new_n330_) | (~new_n326_ & new_n330_))) | (new_n329_ & (~\a[2]  ^ (new_n328_ & (~new_n52_ | ~new_n327_)))) | (~new_n329_ & (~\a[2]  | ~new_n328_ | (new_n52_ & new_n327_)) & (\a[2]  | (new_n328_ & (~new_n52_ | ~new_n327_)))));
  assign new_n326_ = \a[2]  ^ ((~new_n55_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[2]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[4]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[3]  | \a[0]  | ~\a[1] ));
  assign new_n327_ = \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] );
  assign new_n328_ = (~\b[3]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[5]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[4]  | \a[0]  | ~\a[1] );
  assign new_n329_ = (~\a[5]  | ((~\b[0]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[1]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )))) ^ ((~\b[1]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[2]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )));
  assign new_n330_ = ((\b[0]  & (\a[3]  | \a[4] ) & (~\a[3]  | ~\a[4] ) & (\a[2]  ^ ~\a[3] )) | (\b[1]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (\a[4]  ^ ~\a[5] )) | ((\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (\a[4]  | \a[5] ) & (~\a[4]  | ~\a[5] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[5]  & \b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ));
  assign new_n331_ = ((\b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] )) | (\a[2]  & (((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] )) | (~\a[2]  & ((((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )) & ((\b[2]  ^ \b[3] ) | (\b[1]  & (\b[0]  | \b[2] ))) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] ) & ~\a[0]  & ~\a[1] ) | (\b[3]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[2]  & ~\a[0]  & \a[1] )))) & ((\b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (~\a[2]  ^ ((((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] )))) | (\a[2]  & (~\b[1]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[0]  | \a[0]  | ~\a[1] ) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\a[0]  | ~\b[0] ) & (~\b[2]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[1]  | \a[0]  | ~\a[1] ) & (~\b[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & ((\b[2]  ^ (\b[0]  | ~\b[1] )) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))));
  assign new_n332_ = \a[2]  ^ ((~\b[6]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[8]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[7]  | \a[0]  | ~\a[1] ) & ((~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n62_ & (~\b[7]  ^ \b[8] )) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )));
  assign new_n333_ = \a[2]  ^ ((~new_n66_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[5]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[7]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[6]  | \a[0]  | ~\a[1] ));
  assign new_n334_ = (new_n292_ | (~new_n293_ & new_n294_)) ^ (new_n291_ ^ (~\a[5]  ^ (new_n290_ & (~new_n55_ | ~new_n287_))));
  assign new_n335_ = \a[2]  ^ (new_n336_ & (~new_n50_ | ~new_n327_));
  assign new_n336_ = (~\b[4]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[6]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[5]  | \a[0]  | ~\a[1] );
  assign new_n337_ = ~new_n293_ ^ new_n294_;
  assign new_n338_ = \a[2]  ^ ((~new_n96_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[9]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[11]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[10]  | \a[0]  | ~\a[1] ));
  assign new_n339_ = (~new_n282_ ^ new_n283_) ^ ((new_n284_ & ~new_n285_) | (((~new_n286_ & new_n295_) | (~new_n289_ & (new_n286_ | ~new_n295_) & (~new_n286_ | new_n295_))) & (~new_n284_ | new_n285_) & (new_n284_ | ~new_n285_)));
  assign new_n340_ = ~new_n341_ & ((~new_n284_ & new_n285_) | (new_n284_ & ~new_n285_) | ((new_n286_ | ~new_n295_) & (new_n289_ | (~new_n286_ & new_n295_) | (new_n286_ & ~new_n295_)))) & ((~new_n284_ ^ new_n285_) | (~new_n286_ & new_n295_) | (~new_n289_ & (new_n286_ | ~new_n295_) & (~new_n286_ | new_n295_)));
  assign new_n341_ = \a[2]  ^ ((~\b[7]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[9]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[8]  | \a[0]  | ~\a[1] ) & (~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n62_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))));
  assign new_n342_ = ~new_n341_ ^ ((~new_n284_ ^ new_n285_) ^ ((~new_n286_ & new_n295_) | (~new_n289_ & (new_n286_ | ~new_n295_) & (~new_n286_ | new_n295_))));
  assign new_n343_ = \a[2]  ^ ((((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n62_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n62_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[8]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[10]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[9]  | \a[0]  | ~\a[1] ));
  assign new_n344_ = ~new_n345_ & (~new_n280_ | ((new_n298_ | (new_n276_ & ~new_n226_) | (~new_n276_ & new_n226_)) & (new_n281_ | (~new_n298_ & (~new_n276_ | new_n226_) & (new_n276_ | ~new_n226_)) | (new_n298_ & (~new_n276_ ^ ~new_n226_))))) & (new_n280_ | (~new_n298_ & (~new_n276_ | new_n226_) & (new_n276_ | ~new_n226_)) | (~new_n281_ & (new_n298_ | (new_n276_ & ~new_n226_) | (~new_n276_ & new_n226_)) & (~new_n298_ | (new_n276_ ^ ~new_n226_))));
  assign new_n345_ = \a[2]  ^ (((new_n92_ ^ \b[11] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[10]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[11]  | \a[0]  | ~\a[1] ));
  assign new_n346_ = ~new_n345_ ^ (new_n280_ ^ ((~new_n298_ & (~new_n276_ | new_n226_) & (new_n276_ | ~new_n226_)) | (~new_n281_ & (new_n298_ | (new_n276_ & ~new_n226_) | (~new_n276_ & new_n226_)) & (~new_n298_ | (new_n276_ ^ ~new_n226_)))));
  assign new_n347_ = \a[2]  ^ (~\b[11]  | ((\a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (new_n92_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))));
  assign new_n348_ = (new_n270_ | (new_n300_ & (new_n272_ | (~new_n275_ & new_n299_)))) ^ (new_n268_ ^ ~new_n301_);
  assign new_n349_ = new_n300_ ^ (new_n272_ | (~new_n275_ & new_n299_));
  assign new_n350_ = ((\a[5]  & (~new_n239_ | (~new_n212_ & (new_n215_ | ~new_n238_))) & (new_n239_ | new_n212_ | (~new_n215_ & new_n238_))) | (((\a[5]  & (new_n215_ | ~new_n238_) & (~new_n215_ | new_n238_)) | (~new_n267_ & (~\a[5]  | (~new_n215_ & new_n238_) | (new_n215_ & ~new_n238_)) & (\a[5]  | (~new_n215_ ^ new_n238_)))) & (~\a[5]  | (new_n239_ & (new_n212_ | (~new_n215_ & new_n238_))) | (~new_n239_ & ~new_n212_ & (new_n215_ | ~new_n238_))) & (\a[5]  | (new_n239_ ^ (new_n212_ | (~new_n215_ & new_n238_)))))) ^ (\a[5]  ^ (new_n266_ ^ (new_n210_ | (new_n239_ & (new_n212_ | (~new_n215_ & new_n238_))))));
  assign new_n351_ = ((\a[5]  & (~new_n215_ | new_n238_) & (new_n215_ | ~new_n238_)) | (~new_n267_ & (~\a[5]  | (new_n215_ & ~new_n238_) | (~new_n215_ & new_n238_)) & (\a[5]  | (new_n215_ ^ ~new_n238_)))) ^ (\a[5]  ^ (new_n239_ ^ (new_n212_ | (~new_n215_ & new_n238_))));
  assign new_n352_ = ~new_n205_ ^ new_n260_;
  assign new_n353_ = (~new_n261_ | ~\a[5] ) & (((~new_n262_ | ~\a[5] ) & ((new_n262_ & \a[5] ) | (~new_n262_ & ~\a[5] ) | ((~new_n263_ | ~\a[5] ) & (new_n265_ | (new_n263_ & \a[5] ) | (~new_n263_ & ~\a[5] ))))) | (~new_n261_ & ~\a[5] ) | (new_n261_ & \a[5] ));
  assign new_n354_ = ((new_n262_ & \a[5] ) | ((~new_n262_ | ~\a[5] ) & (new_n262_ | \a[5] ) & ((new_n263_ & \a[5] ) | (~new_n265_ & (~new_n263_ | ~\a[5] ) & (new_n263_ | \a[5] ))))) ^ (~new_n261_ ^ ~\a[5] );
  assign new_n355_ = ((new_n256_ & \a[5] ) | ((~new_n256_ | ~\a[5] ) & (new_n256_ | \a[5] ) & ((new_n257_ & \a[5] ) | (((new_n258_ & \a[5] ) | (~new_n259_ & (~new_n258_ | ~\a[5] ) & (new_n258_ | \a[5] ))) & (~new_n257_ | ~\a[5] ) & (new_n257_ | \a[5] ))))) ^ (\a[5]  ^ (~new_n255_ ^ new_n199_));
  assign new_n356_ = ((new_n257_ & \a[5] ) | ((~new_n257_ | ~\a[5] ) & (new_n257_ | \a[5] ) & ((new_n258_ & \a[5] ) | (~new_n259_ & (~new_n258_ | ~\a[5] ) & (new_n258_ | \a[5] ))))) ^ (~new_n256_ ^ ~\a[5] );
  assign new_n357_ = (new_n358_ ^ (~new_n364_ ^ ((~new_n302_ | ~\a[5] ) & (new_n39_ | (new_n302_ & \a[5] ) | (~new_n302_ & ~\a[5] ))))) ^ (~new_n360_ ^ (\a[2]  ^ \a[11] ));
  assign new_n358_ = ~new_n359_ ^ ((~\a[20]  | ((~\a[21]  | ~\b[10] ) & (~\b[11]  | (\a[20]  ^ ~\a[21] )))) & (new_n308_ | (\a[20]  & ((\a[21]  & \b[10] ) | (\b[11]  & (~\a[20]  ^ ~\a[21] )))) | (~\a[20]  & (~\a[21]  | ~\b[11] ))));
  assign new_n359_ = (~\a[11]  | (~new_n305_ & new_n306_) | (new_n305_ & ~new_n306_)) & (((~new_n246_ | ~\a[11] ) & (((~new_n178_ | ~\a[11] ) & (new_n243_ | (new_n178_ & \a[11] ) | (~new_n178_ & ~\a[11] ))) | (new_n246_ & \a[11] ) | (~new_n246_ & ~\a[11] ))) | (~\a[11]  & (new_n305_ ^ new_n306_)) | (\a[11]  & (new_n305_ | ~new_n306_) & (~new_n305_ | new_n306_)));
  assign new_n360_ = new_n361_ ^ (~new_n362_ ^ (~new_n363_ ^ ((~new_n304_ | ~\a[8] ) & ((new_n304_ & \a[8] ) | (~new_n304_ & ~\a[8] ) | ((~new_n303_ | ~\a[8] ) & (new_n40_ | ~new_n242_))))));
  assign new_n361_ = (~new_n307_ | ~\a[17] ) & ((~new_n307_ & ~\a[17] ) | (new_n307_ & \a[17] ) | ((~new_n248_ | ~\a[17] ) & ((new_n248_ & \a[17] ) | (~new_n248_ & ~\a[17] ) | ((~new_n190_ | ~\a[17] ) & ((new_n190_ & \a[17] ) | (~new_n190_ & ~\a[17] ) | ((~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (new_n189_ | (\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~\a[17]  & (new_n194_ ^ new_n186_)))))))));
  assign new_n362_ = ~\a[5]  ^ \a[14] ;
  assign new_n363_ = \a[20]  & (~\a[21]  | ~\b[11] );
  assign new_n364_ = \a[8]  ^ (~\a[17]  ^ ((new_n365_ & \a[14] ) | (~new_n305_ & (new_n365_ | \a[14] ) & (~new_n365_ | ~\a[14] ))));
  assign new_n365_ = (~new_n307_ ^ ~\a[17] ) ^ ((new_n248_ & \a[17] ) | ((~new_n248_ | ~\a[17] ) & (new_n248_ | \a[17] ) & ((new_n190_ & \a[17] ) | ((~new_n190_ | ~\a[17] ) & (new_n190_ | \a[17] ) & ((\a[17]  & (new_n194_ | ~new_n186_) & (~new_n194_ | new_n186_)) | (~new_n189_ & (~\a[17]  | (~new_n194_ & new_n186_) | (new_n194_ & ~new_n186_)) & (\a[17]  | (~new_n194_ ^ new_n186_))))))));
  assign new_n366_ = (((~new_n355_ | ~\a[2] ) & ((new_n355_ & \a[2] ) | (~new_n355_ & ~\a[2] ) | ((~new_n356_ | ~\a[2] ) & (new_n311_ | (new_n356_ & \a[2] ) | (~new_n356_ & ~\a[2] ))))) ^ (\a[2]  ^ (new_n310_ ^ ~new_n254_))) & ((~new_n355_ ^ \a[2] ) ^ ((new_n356_ & \a[2] ) | (~new_n311_ & (~new_n356_ | ~\a[2] ) & (new_n356_ | \a[2] )))) & (new_n311_ ^ (new_n356_ ^ \a[2] )) & ~new_n367_ & new_n368_;
  assign new_n367_ = ((\a[2]  & ((new_n258_ & \a[5] ) | (~new_n258_ & ~\a[5] ) | ((~new_n352_ | ~\a[5] ) & (new_n353_ | (new_n352_ & \a[5] ) | (~new_n352_ & ~\a[5] )))) & ((new_n258_ ^ \a[5] ) | (new_n352_ & \a[5] ) | (~new_n353_ & (~new_n352_ | ~\a[5] ) & (new_n352_ | \a[5] )))) | (((\a[2]  & (new_n353_ | (new_n352_ & \a[5] ) | (~new_n352_ & ~\a[5] )) & (~new_n353_ | (new_n352_ ^ \a[5] ))) | (((new_n354_ & \a[2] ) | (~new_n312_ & (~new_n354_ | ~\a[2] ) & (new_n354_ | \a[2] ))) & (~\a[2]  | (~new_n353_ & (~new_n352_ | ~\a[5] ) & (new_n352_ | \a[5] )) | (new_n353_ & (~new_n352_ ^ \a[5] ))) & (\a[2]  | (~new_n353_ ^ (new_n352_ ^ \a[5] ))))) & (~\a[2]  | ((~new_n258_ | ~\a[5] ) & (new_n258_ | \a[5] ) & ((new_n352_ & \a[5] ) | (~new_n353_ & (~new_n352_ | ~\a[5] ) & (new_n352_ | \a[5] )))) | ((~new_n258_ ^ \a[5] ) & (~new_n352_ | ~\a[5] ) & (new_n353_ | (new_n352_ & \a[5] ) | (~new_n352_ & ~\a[5] )))) & (\a[2]  | ((new_n258_ ^ \a[5] ) ^ ((new_n352_ & \a[5] ) | (~new_n353_ & (~new_n352_ | ~\a[5] ) & (new_n352_ | \a[5] ))))))) ^ (\a[2]  ^ ((new_n257_ ^ \a[5] ) ^ ((new_n258_ & \a[5] ) | ((~new_n258_ | ~\a[5] ) & (new_n258_ | \a[5] ) & ((new_n352_ & \a[5] ) | (~new_n353_ & (~new_n352_ | ~\a[5] ) & (new_n352_ | \a[5] )))))));
  assign new_n368_ = ((~\a[2]  ^ (new_n369_ ^ ~new_n259_)) ^ ((new_n370_ & \a[2] ) | ((~new_n370_ | ~\a[2] ) & (new_n370_ | \a[2] ) & ((new_n354_ & \a[2] ) | ((~new_n354_ | ~\a[2] ) & (new_n354_ | \a[2] ) & ((new_n314_ & \a[2] ) | (~new_n371_ & (~new_n314_ | ~\a[2] ) & (new_n314_ | \a[2] )))))))) & ((~new_n370_ ^ \a[2] ) ^ ((new_n354_ & \a[2] ) | ((~new_n354_ | ~\a[2] ) & (new_n354_ | \a[2] ) & ((new_n314_ & \a[2] ) | (~new_n371_ & (~new_n314_ | ~\a[2] ) & (new_n314_ | \a[2] )))))) & ((new_n354_ ^ \a[2] ) | (new_n314_ & \a[2] ) | (~new_n371_ & (~new_n314_ | ~\a[2] ) & (new_n314_ | \a[2] ))) & ((new_n354_ & \a[2] ) | (~new_n354_ & ~\a[2] ) | ((~new_n314_ | ~\a[2] ) & (new_n371_ | (new_n314_ & \a[2] ) | (~new_n314_ & ~\a[2] )))) & (~new_n371_ | (new_n314_ ^ \a[2] )) & new_n372_ & (new_n371_ | (new_n314_ & \a[2] ) | (~new_n314_ & ~\a[2] ));
  assign new_n369_ = ~new_n258_ ^ ~\a[5] ;
  assign new_n370_ = ~new_n353_ ^ (~new_n352_ ^ ~\a[5] );
  assign new_n371_ = (~\a[2]  | (new_n313_ & ~new_n265_) | (~new_n313_ & new_n265_)) & (((~new_n350_ | ~\a[2] ) & (((~new_n351_ | ~\a[2] ) & (new_n315_ | (new_n351_ & \a[2] ) | (~new_n351_ & ~\a[2] ))) | (new_n350_ & \a[2] ) | (~new_n350_ & ~\a[2] ))) | (\a[2]  & (~new_n313_ | new_n265_) & (new_n313_ | ~new_n265_)) | (~\a[2]  & (~new_n313_ ^ ~new_n265_)));
  assign new_n372_ = ((new_n350_ & \a[2] ) | (((new_n351_ & \a[2] ) | ((~new_n351_ | ~\a[2] ) & (new_n351_ | \a[2] ) & ((new_n316_ & \a[2] ) | (~new_n373_ & (~new_n316_ | ~\a[2] ) & (new_n316_ | \a[2] ))))) & (~new_n350_ | ~\a[2] ) & (new_n350_ | \a[2] )) | (\a[2]  ^ (~new_n313_ ^ new_n265_))) & (((~new_n350_ | ~\a[2] ) & (((~new_n351_ | ~\a[2] ) & ((new_n351_ & \a[2] ) | (~new_n351_ & ~\a[2] ) | ((~new_n316_ | ~\a[2] ) & (new_n373_ | (new_n316_ & \a[2] ) | (~new_n316_ & ~\a[2] ))))) | (new_n350_ & \a[2] ) | (~new_n350_ & ~\a[2] ))) | (\a[2]  & (new_n313_ | ~new_n265_) & (~new_n313_ | new_n265_)) | (~\a[2]  & (new_n313_ ^ new_n265_))) & (((~new_n351_ | ~\a[2] ) & ((new_n351_ & \a[2] ) | (~new_n351_ & ~\a[2] ) | ((~new_n316_ | ~\a[2] ) & (new_n373_ | (new_n316_ & \a[2] ) | (~new_n316_ & ~\a[2] ))))) ^ (new_n350_ ^ \a[2] )) & ((~new_n351_ ^ \a[2] ) ^ ((new_n316_ & \a[2] ) | (~new_n373_ & (~new_n316_ | ~\a[2] ) & (new_n316_ | \a[2] )))) & (~new_n373_ | (new_n316_ ^ \a[2] )) & new_n374_ & (new_n373_ | (new_n316_ & \a[2] ) | (~new_n316_ & ~\a[2] ));
  assign new_n373_ = (~new_n348_ | ~\a[2] ) & ((~new_n348_ & ~\a[2] ) | (new_n348_ & \a[2] ) | ((~new_n349_ | ~\a[2] ) & (new_n318_ | (~new_n349_ & ~\a[2] ) | (new_n349_ & \a[2] ))));
  assign new_n374_ = ((~new_n348_ ^ \a[2] ) ^ ((\a[2]  & (~new_n300_ | (~new_n272_ & (new_n275_ | ~new_n299_))) & (new_n300_ | new_n272_ | (~new_n275_ & new_n299_))) | ((~\a[2]  | (new_n300_ & (new_n272_ | (~new_n275_ & new_n299_))) | (~new_n300_ & ~new_n272_ & (new_n275_ | ~new_n299_))) & (\a[2]  | (new_n300_ ^ (new_n272_ | (~new_n275_ & new_n299_)))) & ((\a[2]  & (new_n275_ | ~new_n299_) & (~new_n275_ | new_n299_)) | (~new_n375_ & (~\a[2]  | (~new_n275_ & new_n299_) | (new_n275_ & ~new_n299_)) & (\a[2]  | (~new_n275_ ^ new_n299_))))))) & ((~\a[2]  ^ (new_n300_ ^ (new_n272_ | (~new_n275_ & new_n299_)))) ^ ((\a[2]  & (new_n275_ | ~new_n299_) & (~new_n275_ | new_n299_)) | (~new_n375_ & (~\a[2]  | (~new_n275_ & new_n299_) | (new_n275_ & ~new_n299_)) & (\a[2]  | (~new_n275_ ^ new_n299_))))) & new_n376_ & (new_n375_ ^ (\a[2]  ^ (~new_n275_ ^ new_n299_)));
  assign new_n375_ = (~new_n319_ | new_n347_) & ((new_n319_ & ~new_n347_) | (~new_n319_ & new_n347_) | (~new_n344_ & (new_n321_ | ~new_n346_)));
  assign new_n376_ = (new_n380_ | new_n344_ | (new_n346_ & (new_n377_ | (~new_n378_ & ~new_n377_ & ~new_n379_)))) & (~new_n380_ | (~new_n344_ & (~new_n346_ | (~new_n377_ & (new_n378_ | new_n377_ | new_n379_))))) & (new_n346_ | new_n377_ | (~new_n378_ & ~new_n377_ & ~new_n379_)) & (~new_n346_ | (~new_n377_ & (new_n378_ | new_n377_ | new_n379_))) & (~new_n378_ | (~new_n377_ & ~new_n379_)) & new_n381_ & (new_n378_ | new_n377_ | new_n379_);
  assign new_n377_ = ~new_n338_ & (new_n322_ | ~new_n281_) & (~new_n322_ | new_n281_);
  assign new_n378_ = (~new_n339_ | new_n343_) & ((new_n339_ & ~new_n343_) | (~new_n339_ & new_n343_) | (~new_n340_ & (new_n323_ | ~new_n342_)));
  assign new_n379_ = new_n338_ & (new_n322_ ^ new_n281_);
  assign new_n380_ = ~new_n347_ ^ (new_n320_ ^ (new_n278_ | (new_n280_ & ((~new_n298_ & (~new_n276_ | new_n226_) & (new_n276_ | ~new_n226_)) | (~new_n281_ & (new_n298_ | (new_n276_ & ~new_n226_) | (~new_n276_ & new_n226_)) & (~new_n298_ | (new_n276_ ^ ~new_n226_)))))));
  assign new_n381_ = (~new_n383_ ^ (new_n340_ | (~new_n323_ & new_n342_))) & (new_n323_ ^ new_n342_) & ~new_n384_ & ~new_n385_ & ~new_n382_ & new_n386_;
  assign new_n382_ = (new_n333_ | ~new_n334_) & (~new_n333_ | new_n334_) & ((~new_n335_ & new_n337_) | (~new_n325_ & (new_n335_ | ~new_n337_) & (~new_n335_ | new_n337_)));
  assign new_n383_ = ~new_n339_ ^ new_n343_;
  assign new_n384_ = (~new_n332_ ^ (new_n324_ ^ ~new_n289_)) ^ ((~new_n333_ & new_n334_) | ((new_n333_ | ~new_n334_) & (~new_n333_ | new_n334_) & ((~new_n335_ & new_n337_) | (~new_n325_ & (new_n335_ | ~new_n337_) & (~new_n335_ | new_n337_)))));
  assign new_n385_ = (new_n333_ ^ new_n334_) & (new_n335_ | ~new_n337_) & (new_n325_ | (~new_n335_ & new_n337_) | (new_n335_ & ~new_n337_));
  assign new_n386_ = (~new_n325_ | new_n387_) & (new_n325_ | ~new_n387_) & (new_n396_ | (~new_n326_ & new_n330_) | (new_n331_ & (new_n326_ | ~new_n330_) & (~new_n326_ | new_n330_))) & (~new_n396_ | ((new_n326_ | ~new_n330_) & (~new_n331_ | (~new_n326_ & new_n330_) | (new_n326_ & ~new_n330_)))) & (~new_n331_ ^ (~new_n326_ ^ new_n330_)) & new_n388_ & ~new_n397_;
  assign new_n387_ = ~new_n335_ ^ new_n337_;
  assign new_n388_ = new_n389_ & (\a[2]  ? (((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[1]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[0]  | \a[0]  | ~\a[1] )) : ((\b[2]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[1]  & ~\a[0]  & \a[1] ) | (\b[0]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | ((~\b[2]  ^ (\b[0]  | ~\b[1] )) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] ))));
  assign new_n389_ = ~new_n390_ & (~new_n391_ | ~new_n392_ | ~new_n393_) & \a[0]  & \b[0]  & (~new_n394_ | ~new_n395_);
  assign new_n390_ = ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[1]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[0]  | \a[0]  | ~\a[1] ) & ((\b[2]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[1]  & ~\a[0]  & \a[1] ) | (\b[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] ) & ~\a[0]  & ~\a[1] ) | (\a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] ) & (~\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n391_ = ~\a[1]  & ~\a[2]  & ~\a[3]  & ~\a[4]  & ~\a[7]  & ~\a[8] ;
  assign new_n392_ = ~\a[13]  & ~\a[14]  & ~\a[11]  & ~\a[12]  & ~\a[5]  & ~\a[6]  & ~\a[9]  & ~\a[10] ;
  assign new_n393_ = ~\a[17]  & ~\a[18]  & ~\a[19]  & ~\a[20]  & ~\a[21]  & ~\a[15]  & ~\a[16] ;
  assign new_n394_ = ~\b[11]  & ~\b[1]  & ~\b[2] ;
  assign new_n395_ = ~\b[9]  & ~\b[10]  & ~\b[7]  & ~\b[8]  & ~\b[3]  & ~\b[4]  & ~\b[5]  & ~\b[6] ;
  assign new_n396_ = new_n329_ ^ (~\a[2]  ^ (new_n328_ & (~new_n52_ | ~new_n327_)));
  assign new_n397_ = (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) ^ (\a[2]  ^ ((((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] )));
  assign new_n398_ = ((new_n250_ & \a[5] ) | ((~new_n250_ | ~\a[5] ) & (new_n250_ | \a[5] ) & ((new_n251_ & \a[5] ) | (((new_n253_ & \a[5] ) | (~new_n254_ & (~new_n253_ | ~\a[5] ) & (new_n253_ | \a[5] ))) & (~new_n251_ | ~\a[5] ) & (new_n251_ | \a[5] ))))) ^ (\a[5]  ^ (~new_n40_ ^ new_n242_));
  assign new_n399_ = ((new_n251_ & \a[5] ) | ((~new_n251_ | ~\a[5] ) & (new_n251_ | \a[5] ) & ((new_n253_ & \a[5] ) | (~new_n254_ & (~new_n253_ | ~\a[5] ) & (new_n253_ | \a[5] ))))) ^ (~new_n250_ ^ ~\a[5] );
  assign new_n400_ = (~new_n251_ ^ ~\a[5] ) ^ ((new_n253_ & \a[5] ) | (~new_n254_ & (new_n253_ | \a[5] ) & (~new_n253_ | ~\a[5] )));
endmodule


