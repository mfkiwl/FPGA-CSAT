// Benchmark "multiplier_448338251_sat" written by ABC on Fri Nov 11 15:31:14 2022

module multiplier_448338251_sat ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] ,
    sat  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] ;
  output sat;
  wire new_n47_, new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_,
    new_n54_, new_n55_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_,
    new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_,
    new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n74_,
    new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_,
    new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_,
    new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_,
    new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_;
  assign sat = (new_n47_ | (~new_n637_ ^ ((new_n525_ & \a[2] ) | (~new_n527_ & (~new_n525_ | ~\a[2] ) & (new_n525_ | \a[2] ))))) & (~new_n47_ | (~new_n637_ & ((new_n525_ & \a[2] ) | (~new_n527_ & (~new_n525_ | ~\a[2] ) & (new_n525_ | \a[2] )))) | (new_n637_ & (~new_n525_ | ~\a[2] ) & (new_n527_ | (new_n525_ & \a[2] ) | (~new_n525_ & ~\a[2] )))) & new_n589_ & (new_n527_ ^ (new_n525_ ^ \a[2] ));
  assign new_n47_ = new_n524_ ^ (new_n48_ ^ (~new_n523_ ^ (~\a[26]  | (\a[27]  & \b[14] ))));
  assign new_n48_ = \a[2]  ^ ((\a[5]  & (~new_n427_ | ((~new_n522_ | ~\a[8] ) & (new_n49_ | (new_n522_ & \a[8] ) | (~new_n522_ & ~\a[8] )))) & (new_n427_ | (new_n522_ & \a[8] ) | (~new_n49_ & (~new_n522_ | ~\a[8] ) & (new_n522_ | \a[8] )))) | (((\a[5]  & (new_n49_ | (new_n522_ & \a[8] ) | (~new_n522_ & ~\a[8] )) & (~new_n49_ | (new_n522_ ^ \a[8] ))) | (((new_n451_ & \a[5] ) | (~new_n452_ & (~new_n451_ | ~\a[5] ) & (new_n451_ | \a[5] ))) & (~\a[5]  | (~new_n49_ & (~new_n522_ | ~\a[8] ) & (new_n522_ | \a[8] )) | (new_n49_ & (~new_n522_ ^ \a[8] ))) & (\a[5]  | (~new_n49_ ^ (new_n522_ ^ \a[8] ))))) & (~\a[5]  | (new_n427_ & ((new_n522_ & \a[8] ) | (~new_n49_ & (~new_n522_ | ~\a[8] ) & (new_n522_ | \a[8] )))) | (~new_n427_ & (~new_n522_ | ~\a[8] ) & (new_n49_ | (new_n522_ & \a[8] ) | (~new_n522_ & ~\a[8] )))) & (\a[5]  | (new_n427_ ^ ((new_n522_ & \a[8] ) | (~new_n49_ & (~new_n522_ | ~\a[8] ) & (new_n522_ | \a[8] )))))));
  assign new_n49_ = (~\a[8]  | ((~new_n379_ | ~\a[11] ) & (new_n379_ | \a[11] ) & ((new_n423_ & \a[11] ) | ((~new_n423_ | ~\a[11] ) & (new_n423_ | \a[11] ) & ((new_n424_ & \a[11] ) | ((~new_n424_ | ~\a[11] ) & (new_n424_ | \a[11] ) & ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] )))))))) | ((~new_n379_ ^ \a[11] ) & (~new_n423_ | ~\a[11] ) & ((new_n423_ & \a[11] ) | (~new_n423_ & ~\a[11] ) | ((~new_n424_ | ~\a[11] ) & ((new_n424_ & \a[11] ) | (~new_n424_ & ~\a[11] ) | ((~new_n425_ | ~\a[11] ) & (new_n426_ | (new_n425_ & \a[11] ) | (~new_n425_ & ~\a[11] )))))))) & (((~\a[8]  | ((~new_n423_ | ~\a[11] ) & (new_n423_ | \a[11] ) & ((new_n424_ & \a[11] ) | ((~new_n424_ | ~\a[11] ) & (new_n424_ | \a[11] ) & ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] )))))) | ((~new_n423_ ^ \a[11] ) & (~new_n424_ | ~\a[11] ) & ((new_n424_ & \a[11] ) | (~new_n424_ & ~\a[11] ) | ((~new_n425_ | ~\a[11] ) & (new_n426_ | (new_n425_ & \a[11] ) | (~new_n425_ & ~\a[11] )))))) & ((\a[8]  & ((new_n423_ & \a[11] ) | (~new_n423_ & ~\a[11] ) | ((~new_n424_ | ~\a[11] ) & ((new_n424_ & \a[11] ) | (~new_n424_ & ~\a[11] ) | ((~new_n425_ | ~\a[11] ) & (new_n426_ | (new_n425_ & \a[11] ) | (~new_n425_ & ~\a[11] )))))) & ((new_n423_ ^ \a[11] ) | (new_n424_ & \a[11] ) | ((~new_n424_ | ~\a[11] ) & (new_n424_ | \a[11] ) & ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] )))))) | (~\a[8]  & ((~new_n423_ ^ \a[11] ) ^ ((new_n424_ & \a[11] ) | ((~new_n424_ | ~\a[11] ) & (new_n424_ | \a[11] ) & ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] ))))))) | ((~\a[8]  | ((~new_n424_ | ~\a[11] ) & (new_n424_ | \a[11] ) & ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] )))) | ((~new_n424_ ^ \a[11] ) & (~new_n425_ | ~\a[11] ) & (new_n426_ | (new_n425_ & \a[11] ) | (~new_n425_ & ~\a[11] )))) & ((\a[8]  & ((new_n424_ & \a[11] ) | (~new_n424_ & ~\a[11] ) | ((~new_n425_ | ~\a[11] ) & (new_n426_ | (new_n425_ & \a[11] ) | (~new_n425_ & ~\a[11] )))) & ((new_n424_ ^ \a[11] ) | (new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] )))) | (~\a[8]  & ((~new_n424_ ^ \a[11] ) ^ ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] ))))) | ((~\a[8]  | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] )) | (new_n426_ & (~new_n425_ ^ \a[11] ))) & (new_n50_ | (\a[8]  & (new_n426_ | (new_n425_ & \a[11] ) | (~new_n425_ & ~\a[11] )) & (~new_n426_ | (new_n425_ ^ \a[11] ))) | (~\a[8]  & (new_n426_ ^ (new_n425_ ^ \a[11] ))))))))) | (\a[8]  & ((new_n379_ & \a[11] ) | (~new_n379_ & ~\a[11] ) | ((~new_n423_ | ~\a[11] ) & ((new_n423_ & \a[11] ) | (~new_n423_ & ~\a[11] ) | ((~new_n424_ | ~\a[11] ) & ((new_n424_ & \a[11] ) | (~new_n424_ & ~\a[11] ) | ((~new_n425_ | ~\a[11] ) & (new_n426_ | (new_n425_ & \a[11] ) | (~new_n425_ & ~\a[11] )))))))) & ((new_n379_ ^ \a[11] ) | (new_n423_ & \a[11] ) | ((~new_n423_ | ~\a[11] ) & (new_n423_ | \a[11] ) & ((new_n424_ & \a[11] ) | ((~new_n424_ | ~\a[11] ) & (new_n424_ | \a[11] ) & ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] )))))))) | (~\a[8]  & ((~new_n379_ ^ \a[11] ) ^ ((new_n423_ & \a[11] ) | ((~new_n423_ | ~\a[11] ) & (new_n423_ | \a[11] ) & ((new_n424_ & \a[11] ) | ((~new_n424_ | ~\a[11] ) & (new_n424_ | \a[11] ) & ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] ))))))))));
  assign new_n50_ = (~new_n51_ | ~\a[8] ) & ((~new_n321_ & (new_n322_ | ~new_n378_)) | (new_n51_ & \a[8] ) | (~new_n51_ & ~\a[8] ));
  assign new_n51_ = (new_n52_ ^ \a[11] ) ^ ((new_n269_ & \a[11] ) | ((~new_n269_ | ~\a[11] ) & (new_n269_ | \a[11] ) & ((\a[11]  & (~new_n270_ | new_n320_) & (new_n270_ | ~new_n320_)) | (~new_n271_ & (~\a[11]  | (new_n270_ & ~new_n320_) | (~new_n270_ & new_n320_)) & (\a[11]  | (new_n270_ ^ ~new_n320_))))));
  assign new_n52_ = (new_n153_ ^ \a[14] ) ^ ((new_n221_ & \a[14] ) | ((~new_n221_ | ~\a[14] ) & (new_n221_ | \a[14] ) & ((\a[14]  & (~new_n53_ | (~new_n176_ & (new_n177_ | ~new_n220_))) & (new_n53_ | new_n176_ | (~new_n177_ & new_n220_))) | (((\a[14]  & (new_n177_ | ~new_n220_) & (~new_n177_ | new_n220_)) | (~new_n222_ & (~\a[14]  | (~new_n177_ & new_n220_) | (new_n177_ & ~new_n220_)) & (\a[14]  | (~new_n177_ ^ new_n220_)))) & (~\a[14]  | (new_n53_ & (new_n176_ | (~new_n177_ & new_n220_))) | (~new_n53_ & ~new_n176_ & (new_n177_ | ~new_n220_))) & (\a[14]  | (new_n53_ ^ (new_n176_ | (~new_n177_ & new_n220_))))))));
  assign new_n53_ = ~new_n54_ ^ ~\a[17] ;
  assign new_n54_ = (new_n115_ | (~new_n118_ & new_n151_)) ^ (~new_n55_ & ~new_n152_);
  assign new_n55_ = ~new_n113_ & (~new_n99_ | ((~new_n110_ | new_n111_) & (new_n56_ | (~new_n110_ & new_n111_) | (new_n110_ & ~new_n111_)))) & (new_n99_ | (new_n110_ & ~new_n111_) | (~new_n56_ & (new_n110_ | ~new_n111_) & (~new_n110_ | new_n111_)));
  assign new_n56_ = (~new_n57_ | new_n96_) & (((~new_n77_ | new_n98_) & ((~new_n78_ & (new_n81_ | ~new_n95_)) | (new_n77_ & ~new_n98_) | (~new_n77_ & new_n98_))) | (new_n57_ & ~new_n96_) | (~new_n57_ & new_n96_));
  assign new_n57_ = new_n74_ ^ (new_n58_ | (new_n73_ & (new_n62_ | (~new_n65_ & new_n72_))));
  assign new_n58_ = ((\b[3]  & (~\a[26]  ^ ~\a[27] )) | (\b[2]  & \a[27]  & (~\a[26]  | \a[27] ) & (\a[26]  | ~\a[27] ))) & (~\a[26]  ^ (new_n61_ & (~new_n59_ | ~new_n60_)));
  assign new_n59_ = (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] ) & (\a[25]  | \a[26] ) & (~\a[25]  | ~\a[26] );
  assign new_n60_ = ((\b[4]  & \b[5] ) | (((\b[3]  & \b[4] ) | (((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))) & (~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ))) & (~\b[4]  | ~\b[5] ) & (\b[4]  | \b[5] ))) ^ (\b[5]  ^ \b[6] );
  assign new_n61_ = (~\b[4]  | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  ^ ~\a[25] )) & (~\b[5]  | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] )) & (~\b[6]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  ^ ~\a[26] ));
  assign new_n62_ = ((\b[2]  & (~\a[26]  ^ ~\a[27] )) | (\b[1]  & \a[27]  & (~\a[26]  | \a[27] ) & (\a[26]  | ~\a[27] ))) & (~\a[26]  ^ (new_n64_ & (~new_n59_ | ~new_n63_)));
  assign new_n63_ = ((\b[3]  & \b[4] ) | (((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))) & (~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ))) ^ (\b[4]  ^ \b[5] );
  assign new_n64_ = (~\b[3]  | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  ^ ~\a[25] )) & (~\b[4]  | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] )) & (~\b[5]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  ^ ~\a[26] ));
  assign new_n65_ = (new_n68_ | (\a[26]  ^ (new_n67_ & (~new_n59_ | ~new_n66_)))) & ((~new_n69_ & (new_n70_ | ~new_n71_)) | (~new_n68_ & (~\a[26]  ^ (new_n67_ & (~new_n59_ | ~new_n66_)))) | (new_n68_ & (~\a[26]  | ~new_n67_ | (new_n59_ & new_n66_)) & (\a[26]  | (new_n67_ & (~new_n59_ | ~new_n66_)))));
  assign new_n66_ = ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))) ^ (\b[3]  ^ \b[4] );
  assign new_n67_ = (~\b[2]  | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  ^ ~\a[25] )) & (~\b[3]  | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] )) & (~\b[4]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  ^ ~\a[26] ));
  assign new_n68_ = (~\b[0]  | ~\a[27]  | (\a[26]  & ~\a[27] ) | (~\a[26]  & \a[27] )) & (~\b[1]  | (\a[26]  ^ ~\a[27] ));
  assign new_n69_ = \b[0]  & (~\a[26]  ^ ~\a[27] ) & (~\b[0]  | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] )) & (~\b[1]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  ^ ~\a[26] )) & ((~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[26]  & (~\b[0]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~\b[0]  | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  ^ ~\a[25] )) & ((~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  ^ ~\a[26] )) & (~\b[1]  | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] ));
  assign new_n70_ = \a[26]  ^ (((~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  ^ ~\a[25] )) & (~\b[3]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  ^ ~\a[26] )) & (~\b[2]  | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] )));
  assign new_n71_ = (\b[0]  & (~\a[26]  ^ ~\a[27] )) ^ ((~\b[0]  | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] )) & (~\b[1]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  ^ ~\a[26] )) & ((~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[26]  & (~\b[0]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~\b[0]  | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  ^ ~\a[25] )) & ((~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  ^ ~\a[26] )) & (~\b[1]  | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] )));
  assign new_n72_ = ((\b[2]  & (~\a[26]  ^ ~\a[27] )) | (\b[1]  & \a[27]  & (~\a[26]  | \a[27] ) & (\a[26]  | ~\a[27] ))) ^ (~\a[26]  ^ (new_n64_ & (~new_n59_ | ~new_n63_)));
  assign new_n73_ = ((\b[3]  & (~\a[26]  ^ ~\a[27] )) | (\b[2]  & \a[27]  & (~\a[26]  | \a[27] ) & (\a[26]  | ~\a[27] ))) ^ (~\a[26]  ^ (new_n61_ & (~new_n59_ | ~new_n60_)));
  assign new_n74_ = ((\b[4]  & (~\a[26]  ^ ~\a[27] )) | (\b[3]  & \a[27]  & (~\a[26]  | \a[27] ) & (\a[26]  | ~\a[27] ))) ^ (~\a[26]  ^ (new_n76_ & (~new_n59_ | ~new_n75_)));
  assign new_n75_ = (\b[6]  ^ \b[7] ) ^ ((\b[5]  & \b[6] ) | (((\b[4]  & \b[5] ) | (((\b[3]  & \b[4] ) | (((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))) & (~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ))) & (~\b[4]  | ~\b[5] ) & (\b[4]  | \b[5] ))) & (~\b[5]  | ~\b[6] ) & (\b[5]  | \b[6] )));
  assign new_n76_ = (~\b[5]  | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  ^ ~\a[25] )) & (~\b[6]  | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] )) & (~\b[7]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  ^ ~\a[26] ));
  assign new_n77_ = new_n73_ ^ (new_n62_ | (~new_n65_ & new_n72_));
  assign new_n78_ = ~new_n79_ & (~new_n65_ | new_n72_) & (new_n65_ | ~new_n72_);
  assign new_n79_ = \a[23]  ^ (((~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n80_ & (~\b[7]  ^ \b[8] )) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~\b[6]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[21]  ^ ~\a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[7]  | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[8]  | (\a[22]  ^ \a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )));
  assign new_n80_ = (~\b[6]  | ~\b[7] ) & ((\b[6]  & \b[7] ) | (~\b[6]  & ~\b[7] ) | ((~\b[5]  | ~\b[6] ) & (((~\b[4]  | ~\b[5] ) & (((~\b[3]  | ~\b[4] ) & (((~\b[2]  | ~\b[3] ) & ((~\b[2]  & ~\b[3] ) | (\b[2]  & \b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] ))) | (\b[3]  & \b[4] ) | (~\b[3]  & ~\b[4] ))) | (\b[4]  & \b[5] ) | (~\b[4]  & ~\b[5] ))) | (\b[5]  & \b[6] ) | (~\b[5]  & ~\b[6] ))));
  assign new_n81_ = (new_n82_ | ~new_n83_) & ((new_n82_ & ~new_n83_) | (~new_n82_ & new_n83_) | ((~new_n84_ | new_n85_) & ((~new_n84_ & new_n85_) | (new_n84_ & ~new_n85_) | ((new_n86_ | ~new_n94_) & (new_n87_ | (~new_n86_ & new_n94_) | (new_n86_ & ~new_n94_))))));
  assign new_n82_ = \a[23]  ^ ((~\b[5]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[21]  ^ ~\a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[6]  | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[7]  | (\a[22]  ^ \a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~new_n75_ | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )));
  assign new_n83_ = (new_n69_ | (~new_n70_ & new_n71_)) ^ (~new_n68_ ^ (~\a[26]  ^ (new_n67_ & (~new_n59_ | ~new_n66_))));
  assign new_n84_ = new_n70_ ^ ~new_n71_;
  assign new_n85_ = \a[23]  ^ ((~\b[4]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[21]  ^ ~\a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[5]  | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[6]  | (\a[22]  ^ \a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~new_n60_ | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )));
  assign new_n86_ = \a[23]  ^ ((~\b[3]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[21]  ^ ~\a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[4]  | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[5]  | (\a[22]  ^ \a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~new_n63_ | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )));
  assign new_n87_ = (~new_n90_ | (\a[23]  ^ (new_n89_ & (~new_n66_ | ~new_n88_)))) & ((~new_n91_ & (new_n92_ | ~new_n93_)) | (new_n90_ & (~\a[23]  ^ (new_n89_ & (~new_n66_ | ~new_n88_)))) | (~new_n90_ & (~\a[23]  | ~new_n89_ | (new_n66_ & new_n88_)) & (\a[23]  | (new_n89_ & (~new_n66_ | ~new_n88_)))));
  assign new_n88_ = (\a[20]  | \a[21] ) & (~\a[20]  | ~\a[21] ) & (\a[22]  | \a[23] ) & (~\a[22]  | ~\a[23] );
  assign new_n89_ = (~\b[2]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & (~\b[3]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[4]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] ));
  assign new_n90_ = ((\b[0]  & (\a[23]  ^ ~\a[24] ) & (\a[24]  | \a[25] ) & (~\a[24]  | ~\a[25] )) | (\b[1]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] ) & (\a[25]  ^ ~\a[26] )) | ((\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] ) & (\a[25]  | \a[26] ) & (~\a[25]  | ~\a[26] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[26]  & \b[0]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] ));
  assign new_n91_ = (~\b[0]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[1]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] )) & ((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[23]  & (~\b[0]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~\b[0]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & ((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] )) & (~\b[1]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & \b[0]  & (~\a[23]  | ~\a[24] ) & (\a[23]  | \a[24] );
  assign new_n92_ = \a[23]  ^ (((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & (~\b[3]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] )) & (~\b[2]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )));
  assign new_n93_ = ((~\b[0]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[1]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] )) & ((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[23]  & (~\b[0]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~\b[0]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & ((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] )) & (~\b[1]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ))) ^ (\b[0]  & (~\a[23]  | ~\a[24] ) & (\a[23]  | \a[24] ));
  assign new_n94_ = ((~\b[0]  | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  ^ ~\a[25] )) & (~\b[1]  | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] )) & (~\b[2]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  ^ ~\a[26] )) & ((~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))) ^ (~\a[26]  | ((~\b[0]  | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] )) & (~\b[1]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  ^ ~\a[26] )) & ((~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[26]  & (~\b[0]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ))));
  assign new_n95_ = ~new_n79_ ^ (new_n65_ ^ ~new_n72_);
  assign new_n96_ = \a[23]  ^ (new_n97_ & (~new_n88_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n97_ = (~\b[8]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & (~\b[9]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[10]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] ));
  assign new_n98_ = \a[23]  ^ ((~\b[7]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[21]  ^ ~\a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[8]  | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[9]  | (\a[22]  ^ \a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & ((\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))));
  assign new_n99_ = ~new_n105_ ^ ((new_n100_ | new_n108_) ^ (~new_n107_ ^ ~new_n109_));
  assign new_n100_ = new_n102_ & (new_n101_ | (new_n74_ & (new_n58_ | (new_n73_ & (new_n62_ | (~new_n65_ & new_n72_))))));
  assign new_n101_ = ((\b[4]  & (~\a[26]  ^ ~\a[27] )) | (\b[3]  & \a[27]  & (~\a[26]  | \a[27] ) & (\a[26]  | ~\a[27] ))) & (~\a[26]  ^ (new_n76_ & (~new_n59_ | ~new_n75_)));
  assign new_n102_ = ~new_n103_ ^ (~\a[26]  ^ (new_n104_ & (~new_n59_ | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n80_ & (~\b[7]  ^ \b[8] )))));
  assign new_n103_ = (~\b[4]  | ~\a[27]  | (\a[26]  & ~\a[27] ) | (~\a[26]  & \a[27] )) & (~\b[5]  | (\a[26]  ^ ~\a[27] ));
  assign new_n104_ = (~\b[6]  | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  ^ ~\a[25] )) & (~\b[7]  | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] )) & (~\b[8]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  ^ ~\a[26] ));
  assign new_n105_ = \a[23]  ^ ((~\b[10]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[21]  ^ ~\a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[11]  | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[12]  | (\a[22]  ^ \a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~new_n106_ | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )));
  assign new_n106_ = (\b[11]  ^ \b[12] ) ^ ((\b[10]  & \b[11] ) | ((~\b[10]  | ~\b[11] ) & (\b[10]  | \b[11] ) & ((\b[9]  & \b[10] ) | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((\b[8]  | \b[9] ) & (~\b[8]  | ~\b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (\b[7]  | \b[8] ) & (~\b[7]  | ~\b[8] )))))))));
  assign new_n107_ = \a[26]  ^ ((~\b[7]  | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (~\a[24]  ^ ~\a[25] ) | (~\a[23]  ^ ~\a[24] )) & (~\b[8]  | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] ) | (~\a[23]  ^ ~\a[24] )) & (~\b[9]  | (\a[25]  ^ \a[26] ) | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & ((\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))));
  assign new_n108_ = ~new_n103_ & (~\a[26]  ^ (new_n104_ & (~new_n59_ | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n80_ & (~\b[7]  ^ \b[8] )))));
  assign new_n109_ = (~\b[5]  | ~\a[27]  | (\a[26]  & ~\a[27] ) | (~\a[26]  & \a[27] )) & (~\b[6]  | (\a[26]  ^ ~\a[27] ));
  assign new_n110_ = new_n102_ ^ (new_n101_ | (new_n74_ & (new_n58_ | (new_n73_ & (new_n62_ | (~new_n65_ & new_n72_))))));
  assign new_n111_ = \a[23]  ^ ((~\b[9]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[21]  ^ ~\a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[10]  | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[11]  | (\a[22]  ^ \a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~new_n112_ | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )));
  assign new_n112_ = (\b[10]  ^ \b[11] ) ^ ((\b[9]  & \b[10] ) | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((\b[8]  | \b[9] ) & (~\b[8]  | ~\b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (\b[7]  | \b[8] ) & (~\b[7]  | ~\b[8] )))))));
  assign new_n113_ = \a[20]  ^ (((\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\b[14]  ^ ((\b[13]  & \b[14] ) | (~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] ))))) & (~\b[14]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[13]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  ^ ~\a[19] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n114_ = (~\b[12]  | ~\b[13] ) & ((\b[12]  & \b[13] ) | (~\b[12]  & ~\b[13] ) | ((~\b[11]  | ~\b[12] ) & ((\b[11]  & \b[12] ) | (~\b[11]  & ~\b[12] ) | ((~\b[10]  | ~\b[11] ) & ((\b[10]  & \b[11] ) | (~\b[10]  & ~\b[11] ) | ((~\b[9]  | ~\b[10] ) & ((\b[9]  & \b[10] ) | (~\b[9]  & ~\b[10] ) | ((~\b[8]  | ~\b[9] ) & ((~\b[8]  & ~\b[9] ) | (\b[8]  & \b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n80_ | (~\b[7]  & ~\b[8] ) | (\b[7]  & \b[8] ))))))))))));
  assign new_n115_ = ~new_n117_ & (~new_n56_ | new_n116_) & (new_n56_ | ~new_n116_);
  assign new_n116_ = new_n110_ ^ ~new_n111_;
  assign new_n117_ = \a[20]  ^ (((~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n114_ & (~\b[13]  ^ \b[14] )) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[13]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[14]  | (\a[19]  ^ \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[12]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  ^ ~\a[19] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n118_ = (~new_n119_ | new_n148_) & ((new_n119_ & ~new_n148_) | (~new_n119_ & new_n148_) | (~new_n121_ & (~new_n147_ | ((~new_n123_ | new_n150_) & (new_n124_ | (new_n123_ & ~new_n150_) | (~new_n123_ & new_n150_))))));
  assign new_n119_ = new_n120_ ^ ((new_n77_ & ~new_n98_) | ((new_n78_ | (~new_n81_ & new_n95_)) & (~new_n77_ | new_n98_) & (new_n77_ | ~new_n98_)));
  assign new_n120_ = ~new_n96_ ^ (new_n74_ ^ (new_n58_ | (new_n73_ & (new_n62_ | (~new_n65_ & new_n72_)))));
  assign new_n121_ = ~new_n122_ & ((~new_n78_ & (new_n81_ | ~new_n95_)) | (new_n77_ & ~new_n98_) | (~new_n77_ & new_n98_)) & (new_n78_ | (~new_n81_ & new_n95_) | (new_n77_ ^ ~new_n98_));
  assign new_n122_ = \a[20]  ^ ((~new_n106_ | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[11]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[12]  | (\a[19]  ^ \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[10]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  ^ ~\a[19] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n123_ = new_n81_ ^ ~new_n95_;
  assign new_n124_ = (~new_n126_ | new_n144_) & ((new_n126_ & ~new_n144_) | (~new_n126_ & new_n144_) | (~new_n127_ & (~new_n143_ | ((new_n146_ | (new_n125_ & ~new_n87_) | (~new_n125_ & new_n87_)) & (new_n129_ | (~new_n146_ & (~new_n125_ | new_n87_) & (new_n125_ | ~new_n87_)) | (new_n146_ & (~new_n125_ ^ ~new_n87_)))))));
  assign new_n125_ = new_n86_ ^ ~new_n94_;
  assign new_n126_ = (new_n82_ ^ ~new_n83_) ^ ((new_n84_ & ~new_n85_) | ((new_n84_ | ~new_n85_) & (~new_n84_ | new_n85_) & ((~new_n86_ & new_n94_) | (~new_n87_ & (new_n86_ | ~new_n94_) & (~new_n86_ | new_n94_)))));
  assign new_n127_ = ~new_n128_ & ((new_n84_ & ~new_n85_) | (~new_n84_ & new_n85_) | ((new_n86_ | ~new_n94_) & (new_n87_ | (~new_n86_ & new_n94_) | (new_n86_ & ~new_n94_)))) & ((new_n84_ ^ ~new_n85_) | (~new_n86_ & new_n94_) | (~new_n87_ & (new_n86_ | ~new_n94_) & (~new_n86_ | new_n94_)));
  assign new_n128_ = \a[20]  ^ (((\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[9]  | (\a[19]  ^ \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[7]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  ^ ~\a[19] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n129_ = (new_n130_ | ~new_n131_) & ((new_n130_ & ~new_n131_) | (~new_n130_ & new_n131_) | ((~new_n132_ | new_n133_) & ((~new_n132_ & new_n133_) | (new_n132_ & ~new_n133_) | ((new_n134_ | ~new_n142_) & (new_n135_ | (~new_n134_ & new_n142_) | (new_n134_ & ~new_n142_))))));
  assign new_n130_ = \a[20]  ^ ((~new_n75_ | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[6]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[7]  | (\a[19]  ^ \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[5]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  ^ ~\a[19] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n131_ = (new_n91_ | (~new_n92_ & new_n93_)) ^ (new_n90_ ^ (~\a[23]  ^ (new_n89_ & (~new_n66_ | ~new_n88_))));
  assign new_n132_ = new_n92_ ^ ~new_n93_;
  assign new_n133_ = \a[20]  ^ ((~new_n60_ | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[5]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[6]  | (\a[19]  ^ \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[4]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  ^ ~\a[19] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n134_ = \a[20]  ^ ((~new_n63_ | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[4]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[5]  | (\a[19]  ^ \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[3]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  ^ ~\a[19] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n135_ = (~new_n138_ | (\a[20]  ^ (new_n137_ & (~new_n66_ | ~new_n136_)))) & ((~new_n139_ & (new_n140_ | ~new_n141_)) | (new_n138_ & (~\a[20]  ^ (new_n137_ & (~new_n66_ | ~new_n136_)))) | (~new_n138_ & (~\a[20]  | ~new_n137_ | (new_n66_ & new_n136_)) & (\a[20]  | (new_n137_ & (~new_n66_ | ~new_n136_)))));
  assign new_n136_ = (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ) & (\a[19]  | \a[20] ) & (~\a[19]  | ~\a[20] );
  assign new_n137_ = (~\b[3]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[4]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & (~\b[2]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ));
  assign new_n138_ = ((\b[0]  & (\a[20]  ^ ~\a[21] ) & (\a[21]  | \a[22] ) & (~\a[21]  | ~\a[22] )) | (\b[1]  & (\a[20]  | \a[21] ) & (~\a[20]  | ~\a[21] ) & (\a[22]  ^ ~\a[23] )) | ((\a[20]  | \a[21] ) & (~\a[20]  | ~\a[21] ) & (\a[22]  | \a[23] ) & (~\a[22]  | ~\a[23] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[23]  & \b[0]  & (\a[20]  | \a[21] ) & (~\a[20]  | ~\a[21] ));
  assign new_n139_ = \b[0]  & (~\a[20]  | ~\a[21] ) & (\a[20]  | \a[21] ) & (~\b[0]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[1]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[20]  & (~\b[0]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & (~\b[1]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[0]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ));
  assign new_n140_ = \a[20]  ^ (((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & (~\b[2]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[1]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] )));
  assign new_n141_ = (\b[0]  & (~\a[20]  | ~\a[21] ) & (\a[20]  | \a[21] )) ^ ((~\b[0]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[1]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[20]  & (~\b[0]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & (~\b[1]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[0]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] )));
  assign new_n142_ = ((~\b[0]  | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  ^ ~\a[22] )) & (~\b[1]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[2]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] )) & ((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))) ^ (~\a[23]  | ((~\b[0]  | (~\a[20]  ^ ~\a[21] ) | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] )) & (~\b[1]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  ^ ~\a[23] )) & ((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\a[22]  & ~\a[23] ) | (\a[22]  & \a[23] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[23]  & (~\b[0]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ))));
  assign new_n143_ = ~new_n128_ ^ ((new_n84_ ^ ~new_n85_) ^ ((~new_n86_ & new_n94_) | (~new_n87_ & (new_n86_ | ~new_n94_) & (~new_n86_ | new_n94_))));
  assign new_n144_ = \a[20]  ^ (new_n145_ & (~new_n136_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n145_ = (~\b[9]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[10]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & (~\b[8]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] ));
  assign new_n146_ = \a[20]  ^ (((~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n80_ & (~\b[7]  ^ \b[8] )) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[7]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[8]  | (\a[19]  ^ \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[6]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  ^ ~\a[19] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n147_ = ~new_n122_ ^ ((new_n78_ | (~new_n81_ & new_n95_)) ^ (new_n77_ ^ ~new_n98_));
  assign new_n148_ = \a[20]  ^ ((~new_n149_ | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[12]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[13]  | (\a[19]  ^ \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[11]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  ^ ~\a[19] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n149_ = (\b[12]  ^ \b[13] ) ^ ((\b[11]  & \b[12] ) | ((~\b[11]  | ~\b[12] ) & (\b[11]  | \b[12] ) & ((\b[10]  & \b[11] ) | ((~\b[10]  | ~\b[11] ) & (\b[10]  | \b[11] ) & ((\b[9]  & \b[10] ) | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((\b[8]  | \b[9] ) & (~\b[8]  | ~\b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (\b[7]  | \b[8] ) & (~\b[7]  | ~\b[8] )))))))))));
  assign new_n150_ = \a[20]  ^ ((~new_n112_ | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[10]  | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] ) | (~\a[17]  ^ ~\a[18] )) & (~\b[11]  | (\a[19]  ^ \a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[9]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  ^ ~\a[19] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n151_ = ~new_n117_ ^ (new_n56_ ^ ~new_n116_);
  assign new_n152_ = new_n113_ & (~new_n99_ ^ ((new_n110_ & ~new_n111_) | (~new_n56_ & (new_n110_ | ~new_n111_) & (~new_n110_ | new_n111_))));
  assign new_n153_ = ((new_n174_ & \a[17] ) | ((~new_n174_ | ~\a[17] ) & (new_n174_ | \a[17] ) & ((new_n54_ & \a[17] ) | ((~new_n54_ | ~\a[17] ) & (new_n54_ | \a[17] ) & (new_n176_ | (~new_n177_ & new_n220_)))))) ^ (\a[17]  ^ (new_n154_ ^ ~new_n165_));
  assign new_n154_ = (~new_n155_ | new_n163_) & ((~new_n55_ & (new_n55_ | new_n152_ | (~new_n115_ & (new_n118_ | ~new_n151_)))) | (new_n155_ & ~new_n163_) | (~new_n155_ & new_n163_));
  assign new_n155_ = new_n157_ ^ (new_n156_ | (new_n99_ & ((new_n110_ & ~new_n111_) | (~new_n56_ & (new_n110_ | ~new_n111_) & (~new_n110_ | new_n111_)))));
  assign new_n156_ = ~new_n105_ & ((~new_n100_ & ~new_n108_) | (~new_n107_ & ~new_n109_) | (new_n107_ & new_n109_)) & (new_n100_ | new_n108_ | (~new_n107_ ^ ~new_n109_));
  assign new_n157_ = ~new_n162_ ^ (new_n158_ ^ ((~new_n107_ & ~new_n109_) | ((new_n100_ | new_n108_) & (new_n107_ | new_n109_) & (~new_n107_ | ~new_n109_))));
  assign new_n158_ = ~new_n161_ ^ (new_n159_ ^ ~\a[26] );
  assign new_n159_ = new_n160_ & (~new_n59_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))))));
  assign new_n160_ = (~\b[8]  | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  ^ ~\a[25] )) & (~\b[9]  | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] )) & (~\b[10]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  ^ ~\a[26] ));
  assign new_n161_ = (~\b[6]  | ~\a[27]  | (\a[26]  & ~\a[27] ) | (~\a[26]  & \a[27] )) & (~\b[7]  | (\a[26]  ^ ~\a[27] ));
  assign new_n162_ = \a[23]  ^ ((~\b[11]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[21]  ^ ~\a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[12]  | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[13]  | (\a[22]  ^ \a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~new_n149_ | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )));
  assign new_n163_ = \a[20]  ^ (~\b[14]  | (((~\a[17]  ^ ~\a[18] ) | (~\a[18]  ^ ~\a[19] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )) & (new_n164_ | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ))));
  assign new_n164_ = (~\b[13]  | ~\b[14] ) & (new_n114_ | (~\b[13]  & ~\b[14] ) | (\b[13]  & \b[14] ));
  assign new_n165_ = ~new_n166_ ^ ~\a[20] ;
  assign new_n166_ = new_n168_ ^ (new_n167_ | (new_n157_ & (new_n156_ | (new_n99_ & ((new_n110_ & ~new_n111_) | (~new_n56_ & (~new_n110_ | new_n111_) & (new_n110_ | ~new_n111_)))))));
  assign new_n167_ = ~new_n162_ & (~new_n158_ | ((new_n107_ | new_n109_) & ((~new_n100_ & ~new_n108_) | (~new_n107_ & ~new_n109_) | (new_n107_ & new_n109_)))) & (new_n158_ | (~new_n107_ & ~new_n109_) | ((new_n100_ | new_n108_) & (new_n107_ | new_n109_) & (~new_n107_ | ~new_n109_)));
  assign new_n168_ = ~new_n173_ ^ (new_n170_ ^ ((~new_n169_ & ~new_n161_) | (((~new_n107_ & ~new_n109_) | ((new_n100_ | new_n108_) & (~new_n107_ | ~new_n109_) & (new_n107_ | new_n109_))) & (new_n169_ | new_n161_) & (~new_n169_ | ~new_n161_))));
  assign new_n169_ = ~new_n159_ ^ ~\a[26] ;
  assign new_n170_ = (new_n171_ ^ ~\a[26] ) ^ ((\b[8]  & (\a[26]  ^ \a[27] )) | (\b[7]  & \a[27]  & (\a[26]  | ~\a[27] ) & (~\a[26]  | \a[27] )));
  assign new_n171_ = new_n172_ & (~new_n59_ | ((~\b[10]  | ~\b[11] ) & (\b[10]  | \b[11] ) & ((\b[9]  & \b[10] ) | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))))) | ((~\b[10]  ^ \b[11] ) & (~\b[9]  | ~\b[10] ) & ((\b[9]  & \b[10] ) | (~\b[9]  & ~\b[10] ) | ((~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))))))));
  assign new_n172_ = (~\b[9]  | (~\a[25]  & ~\a[26] ) | (\a[25]  & \a[26] ) | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  ^ ~\a[25] )) & (~\b[10]  | (~\a[23]  ^ ~\a[24] ) | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] )) & (~\b[11]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\a[25]  ^ ~\a[26] ));
  assign new_n173_ = \a[23]  ^ (((~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n114_ & (~\b[13]  ^ \b[14] )) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~\b[12]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[21]  ^ ~\a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[13]  | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[14]  | (\a[22]  ^ \a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )));
  assign new_n174_ = new_n175_ ^ (new_n55_ | ((new_n115_ | (~new_n118_ & new_n151_)) & ~new_n55_ & ~new_n152_));
  assign new_n175_ = ~new_n163_ ^ (new_n157_ ^ (new_n156_ | (new_n99_ & ((new_n110_ & ~new_n111_) | (~new_n56_ & (new_n110_ | ~new_n111_) & (~new_n110_ | new_n111_))))));
  assign new_n176_ = \a[17]  & (~new_n118_ | new_n151_) & (new_n118_ | ~new_n151_);
  assign new_n177_ = (~new_n178_ | new_n218_) & ((new_n178_ & ~new_n218_) | (~new_n178_ & new_n218_) | (~new_n180_ & (((new_n219_ | (~new_n124_ & new_n217_) | (new_n124_ & ~new_n217_)) & (new_n182_ | (~new_n219_ & (new_n124_ | ~new_n217_) & (~new_n124_ | new_n217_)) | (new_n219_ & (new_n124_ ^ new_n217_)))) | new_n180_ | new_n216_)));
  assign new_n178_ = new_n179_ ^ (new_n121_ | (new_n147_ & ((new_n123_ & ~new_n150_) | (~new_n124_ & (new_n123_ | ~new_n150_) & (~new_n123_ | new_n150_)))));
  assign new_n179_ = ~new_n148_ ^ (new_n120_ ^ ((new_n77_ & ~new_n98_) | ((new_n78_ | (~new_n81_ & new_n95_)) & (~new_n77_ | new_n98_) & (new_n77_ | ~new_n98_))));
  assign new_n180_ = ~new_n181_ & (~new_n147_ | ((~new_n123_ | new_n150_) & (new_n124_ | (new_n123_ & ~new_n150_) | (~new_n123_ & new_n150_)))) & (new_n147_ | (new_n123_ & ~new_n150_) | (~new_n124_ & (~new_n123_ | new_n150_) & (new_n123_ | ~new_n150_)));
  assign new_n181_ = \a[17]  ^ (((\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\b[14]  ^ ((\b[13]  & \b[14] ) | (~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] ))))) & (~\b[14]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[13]  | (~\a[15]  ^ ~\a[16] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n182_ = (~new_n183_ | new_n215_) & ((~new_n185_ & (~new_n214_ | (~new_n187_ & (new_n190_ | ~new_n213_)))) | (new_n183_ & ~new_n215_) | (~new_n183_ & new_n215_));
  assign new_n183_ = new_n184_ ^ (new_n127_ | (new_n143_ & ((~new_n146_ & (new_n87_ | (~new_n86_ & new_n94_) | (new_n86_ & ~new_n94_)) & (~new_n87_ | (~new_n86_ ^ new_n94_))) | (~new_n129_ & (new_n146_ | (~new_n87_ & (new_n86_ | ~new_n94_) & (~new_n86_ | new_n94_)) | (new_n87_ & (new_n86_ ^ new_n94_))) & (~new_n146_ | (~new_n87_ ^ (~new_n86_ ^ new_n94_)))))));
  assign new_n184_ = ~new_n144_ ^ ((new_n82_ ^ ~new_n83_) ^ ((new_n84_ & ~new_n85_) | ((new_n84_ | ~new_n85_) & (~new_n84_ | new_n85_) & ((~new_n86_ & new_n94_) | (~new_n87_ & (new_n86_ | ~new_n94_) & (~new_n86_ | new_n94_))))));
  assign new_n185_ = ~new_n186_ & (~new_n143_ | ((new_n146_ | (~new_n87_ & (new_n86_ | ~new_n94_) & (~new_n86_ | new_n94_)) | (new_n87_ & (new_n86_ ^ new_n94_))) & (new_n129_ | (~new_n146_ & (new_n87_ | (~new_n86_ & new_n94_) | (new_n86_ & ~new_n94_)) & (~new_n87_ | (~new_n86_ ^ new_n94_))) | (new_n146_ & (new_n87_ ^ (~new_n86_ ^ new_n94_)))))) & (new_n143_ | (~new_n146_ & (new_n87_ | (~new_n86_ & new_n94_) | (new_n86_ & ~new_n94_)) & (~new_n87_ | (~new_n86_ ^ new_n94_))) | (~new_n129_ & (new_n146_ | (~new_n87_ & (new_n86_ | ~new_n94_) & (~new_n86_ | new_n94_)) | (new_n87_ & (new_n86_ ^ new_n94_))) & (~new_n146_ | (~new_n87_ ^ (~new_n86_ ^ new_n94_)))));
  assign new_n186_ = \a[17]  ^ ((~new_n106_ | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[11]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[12]  | (\a[16]  ^ \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[10]  | (~\a[15]  ^ ~\a[16] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n187_ = ~new_n189_ & (~new_n129_ | new_n188_) & (new_n129_ | ~new_n188_);
  assign new_n188_ = ~new_n146_ ^ (~new_n87_ ^ (new_n86_ ^ ~new_n94_));
  assign new_n189_ = \a[17]  ^ ((~new_n112_ | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[10]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[11]  | (\a[16]  ^ \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[9]  | (~\a[15]  ^ ~\a[16] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n190_ = (~new_n192_ | new_n210_) & ((new_n192_ & ~new_n210_) | (~new_n192_ & new_n210_) | (~new_n193_ & (~new_n209_ | ((new_n212_ | (new_n191_ & ~new_n135_) | (~new_n191_ & new_n135_)) & (new_n195_ | (~new_n212_ & (~new_n191_ | new_n135_) & (new_n191_ | ~new_n135_)) | (new_n212_ & (~new_n191_ ^ ~new_n135_)))))));
  assign new_n191_ = new_n134_ ^ ~new_n142_;
  assign new_n192_ = (new_n130_ ^ ~new_n131_) ^ ((new_n132_ & ~new_n133_) | ((new_n132_ | ~new_n133_) & (~new_n132_ | new_n133_) & ((~new_n134_ & new_n142_) | (~new_n135_ & (new_n134_ | ~new_n142_) & (~new_n134_ | new_n142_)))));
  assign new_n193_ = ~new_n194_ & ((new_n132_ & ~new_n133_) | (~new_n132_ & new_n133_) | ((new_n134_ | ~new_n142_) & (new_n135_ | (~new_n134_ & new_n142_) | (new_n134_ & ~new_n142_)))) & ((new_n132_ ^ ~new_n133_) | (~new_n134_ & new_n142_) | (~new_n135_ & (new_n134_ | ~new_n142_) & (~new_n134_ | new_n142_)));
  assign new_n194_ = \a[17]  ^ (((\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[9]  | (\a[16]  ^ \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[7]  | (~\a[15]  ^ ~\a[16] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n195_ = (new_n196_ | ~new_n197_) & ((new_n196_ & ~new_n197_) | (~new_n196_ & new_n197_) | ((~new_n198_ | new_n199_) & ((~new_n198_ & new_n199_) | (new_n198_ & ~new_n199_) | ((new_n200_ | ~new_n208_) & (new_n201_ | (~new_n200_ & new_n208_) | (new_n200_ & ~new_n208_))))));
  assign new_n196_ = \a[17]  ^ ((~new_n75_ | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[6]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[7]  | (\a[16]  ^ \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[5]  | (~\a[15]  ^ ~\a[16] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n197_ = (new_n139_ | (~new_n140_ & new_n141_)) ^ (new_n138_ ^ (~\a[20]  ^ (new_n137_ & (~new_n66_ | ~new_n136_))));
  assign new_n198_ = new_n140_ ^ ~new_n141_;
  assign new_n199_ = \a[17]  ^ ((~new_n60_ | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[5]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[6]  | (\a[16]  ^ \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[4]  | (~\a[15]  ^ ~\a[16] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n200_ = \a[17]  ^ ((~new_n63_ | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[4]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[5]  | (\a[16]  ^ \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[3]  | (~\a[15]  ^ ~\a[16] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n201_ = (~new_n204_ | (\a[17]  ^ (new_n203_ & (~new_n66_ | ~new_n202_)))) & ((~new_n205_ & (new_n206_ | ~new_n207_)) | (new_n204_ & (~\a[17]  ^ (new_n203_ & (~new_n66_ | ~new_n202_)))) | (~new_n204_ & (~\a[17]  | ~new_n203_ | (new_n66_ & new_n202_)) & (\a[17]  | (new_n203_ & (~new_n66_ | ~new_n202_)))));
  assign new_n202_ = (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ) & (\a[16]  | \a[17] ) & (~\a[16]  | ~\a[17] );
  assign new_n203_ = (~\b[3]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[4]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & (~\b[2]  | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ));
  assign new_n204_ = ((\b[0]  & (\a[17]  ^ ~\a[18] ) & (\a[18]  | \a[19] ) & (~\a[18]  | ~\a[19] )) | (\b[1]  & (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ) & (\a[19]  ^ ~\a[20] )) | ((\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ) & (\a[19]  | \a[20] ) & (~\a[19]  | ~\a[20] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[20]  & \b[0]  & (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ));
  assign new_n205_ = \b[0]  & (~\a[17]  | ~\a[18] ) & (\a[17]  | \a[18] ) & (~\b[0]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[1]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[17]  & (~\b[0]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & (~\b[1]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[0]  | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ));
  assign new_n206_ = \a[17]  ^ (((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & (~\b[2]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[1]  | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] )));
  assign new_n207_ = (\b[0]  & (~\a[17]  | ~\a[18] ) & (\a[17]  | \a[18] )) ^ ((~\b[0]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[1]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[17]  & (~\b[0]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & (~\b[1]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[0]  | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] )));
  assign new_n208_ = (~\a[20]  | ((~\b[0]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[1]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[20]  & (~\b[0]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )))) ^ ((~\b[1]  | (~\a[17]  ^ ~\a[18] ) | (~\a[18]  & ~\a[19] ) | (\a[18]  & \a[19] )) & (~\b[2]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  ^ ~\a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[17]  ^ ~\a[18] ) | (~\a[19]  & ~\a[20] ) | (\a[19]  & \a[20] ) | (~\a[18]  ^ ~\a[19] )));
  assign new_n209_ = ~new_n194_ ^ ((new_n132_ ^ ~new_n133_) ^ ((~new_n134_ & new_n142_) | (~new_n135_ & (new_n134_ | ~new_n142_) & (~new_n134_ | new_n142_))));
  assign new_n210_ = \a[17]  ^ (new_n211_ & (~new_n202_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n211_ = (~\b[9]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[10]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & (~\b[8]  | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ));
  assign new_n212_ = \a[17]  ^ (((~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n80_ & (~\b[7]  ^ \b[8] )) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[7]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[8]  | (\a[16]  ^ \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[6]  | (~\a[15]  ^ ~\a[16] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n213_ = ~new_n189_ ^ (new_n129_ ^ ~new_n188_);
  assign new_n214_ = ~new_n186_ ^ (new_n143_ ^ ((~new_n146_ & (new_n87_ | (~new_n86_ & new_n94_) | (new_n86_ & ~new_n94_)) & (~new_n87_ | (~new_n86_ ^ new_n94_))) | (~new_n129_ & (new_n146_ | (~new_n87_ & (new_n86_ | ~new_n94_) & (~new_n86_ | new_n94_)) | (new_n87_ & (new_n86_ ^ new_n94_))) & (~new_n146_ | (~new_n87_ ^ (~new_n86_ ^ new_n94_))))));
  assign new_n215_ = \a[17]  ^ ((~new_n149_ | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[12]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[13]  | (\a[16]  ^ \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[11]  | (~\a[15]  ^ ~\a[16] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n216_ = new_n181_ & (~new_n147_ ^ ((~new_n150_ & (new_n81_ | ~new_n95_) & (~new_n81_ | new_n95_)) | (~new_n124_ & (new_n150_ | (~new_n81_ & new_n95_) | (new_n81_ & ~new_n95_)) & (~new_n150_ | (~new_n81_ ^ new_n95_)))));
  assign new_n217_ = ~new_n150_ ^ (new_n81_ ^ ~new_n95_);
  assign new_n218_ = \a[17]  ^ (~\b[14]  | ((new_n164_ | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & ((~\a[15]  ^ ~\a[16] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] ))));
  assign new_n219_ = \a[17]  ^ (((~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n114_ & (~\b[13]  ^ \b[14] )) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[13]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[14]  | (\a[16]  ^ \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[12]  | (~\a[15]  ^ ~\a[16] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n220_ = \a[17]  ^ (new_n118_ ^ ~new_n151_);
  assign new_n221_ = (new_n174_ ^ \a[17] ) ^ ((new_n54_ & \a[17] ) | ((~new_n54_ | ~\a[17] ) & (new_n54_ | \a[17] ) & (new_n176_ | (~new_n177_ & new_n220_))));
  assign new_n222_ = (~new_n223_ | ~\a[14] ) & ((new_n223_ & \a[14] ) | (~new_n223_ & ~\a[14] ) | ((~new_n225_ | ~\a[14] ) & (((~new_n226_ | ~\a[14] ) & (new_n228_ | (~new_n226_ & ~\a[14] ) | (new_n226_ & \a[14] ))) | (new_n225_ & \a[14] ) | (~new_n225_ & ~\a[14] ))));
  assign new_n223_ = new_n224_ ^ (new_n180_ | (~new_n180_ & ~new_n216_ & ((~new_n219_ & (new_n124_ | ~new_n217_) & (~new_n124_ | new_n217_)) | (~new_n182_ & (new_n219_ | (~new_n124_ & new_n217_) | (new_n124_ & ~new_n217_)) & (~new_n219_ | (~new_n124_ ^ new_n217_))))));
  assign new_n224_ = ~new_n218_ ^ (new_n179_ ^ (new_n121_ | (new_n147_ & ((new_n123_ & ~new_n150_) | (~new_n124_ & (~new_n123_ | new_n150_) & (new_n123_ | ~new_n150_))))));
  assign new_n225_ = (~new_n180_ & ~new_n216_) ^ ((~new_n219_ & (~new_n124_ | new_n217_) & (new_n124_ | ~new_n217_)) | (~new_n182_ & (~new_n219_ | (new_n124_ ^ ~new_n217_)) & (new_n219_ | (new_n124_ & ~new_n217_) | (~new_n124_ & new_n217_))));
  assign new_n226_ = new_n182_ ^ ~new_n227_;
  assign new_n227_ = ~new_n219_ ^ (new_n124_ ^ ~new_n217_);
  assign new_n228_ = (~new_n229_ | new_n267_) & ((new_n229_ & ~new_n267_) | (~new_n229_ & new_n267_) | (~new_n230_ & (((new_n268_ | (~new_n190_ & new_n213_) | (new_n190_ & ~new_n213_)) & (new_n232_ | (~new_n268_ & (new_n190_ | ~new_n213_) & (~new_n190_ | new_n213_)) | (new_n268_ & (new_n190_ ^ new_n213_)))) | new_n230_ | new_n266_)));
  assign new_n229_ = (new_n185_ | (new_n214_ & (new_n187_ | (~new_n190_ & new_n213_)))) ^ (new_n183_ ^ ~new_n215_);
  assign new_n230_ = ~new_n231_ & (~new_n214_ | (~new_n187_ & (new_n190_ | ~new_n213_))) & (new_n214_ | new_n187_ | (~new_n190_ & new_n213_));
  assign new_n231_ = \a[14]  ^ (((\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\b[14]  ^ ((\b[13]  & \b[14] ) | (~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] ))))) & (~\b[14]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[13]  | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n232_ = (~new_n233_ | new_n265_) & ((~new_n235_ & (~new_n264_ | (~new_n237_ & (new_n240_ | ~new_n263_)))) | (new_n233_ & ~new_n265_) | (~new_n233_ & new_n265_));
  assign new_n233_ = new_n234_ ^ (new_n193_ | (new_n209_ & ((~new_n212_ & (new_n135_ | (~new_n134_ & new_n142_) | (new_n134_ & ~new_n142_)) & (~new_n135_ | (~new_n134_ ^ new_n142_))) | (~new_n195_ & (new_n212_ | (~new_n135_ & (new_n134_ | ~new_n142_) & (~new_n134_ | new_n142_)) | (new_n135_ & (new_n134_ ^ new_n142_))) & (~new_n212_ | (~new_n135_ ^ (~new_n134_ ^ new_n142_)))))));
  assign new_n234_ = ~new_n210_ ^ ((new_n130_ ^ ~new_n131_) ^ ((new_n132_ & ~new_n133_) | ((new_n132_ | ~new_n133_) & (~new_n132_ | new_n133_) & ((~new_n134_ & new_n142_) | (~new_n135_ & (new_n134_ | ~new_n142_) & (~new_n134_ | new_n142_))))));
  assign new_n235_ = ~new_n236_ & (~new_n209_ | ((new_n212_ | (~new_n135_ & (new_n134_ | ~new_n142_) & (~new_n134_ | new_n142_)) | (new_n135_ & (new_n134_ ^ new_n142_))) & (new_n195_ | (~new_n212_ & (new_n135_ | (~new_n134_ & new_n142_) | (new_n134_ & ~new_n142_)) & (~new_n135_ | (~new_n134_ ^ new_n142_))) | (new_n212_ & (new_n135_ ^ (~new_n134_ ^ new_n142_)))))) & (new_n209_ | (~new_n212_ & (new_n135_ | (~new_n134_ & new_n142_) | (new_n134_ & ~new_n142_)) & (~new_n135_ | (~new_n134_ ^ new_n142_))) | (~new_n195_ & (new_n212_ | (~new_n135_ & (new_n134_ | ~new_n142_) & (~new_n134_ | new_n142_)) | (new_n135_ & (new_n134_ ^ new_n142_))) & (~new_n212_ | (~new_n135_ ^ (~new_n134_ ^ new_n142_)))));
  assign new_n236_ = \a[14]  ^ ((~new_n106_ | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[11]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[12]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[10]  | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n237_ = ~new_n239_ & (~new_n195_ | new_n238_) & (new_n195_ | ~new_n238_);
  assign new_n238_ = ~new_n212_ ^ (~new_n135_ ^ (new_n134_ ^ ~new_n142_));
  assign new_n239_ = \a[14]  ^ ((~new_n112_ | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[10]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[11]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[9]  | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n240_ = (~new_n242_ | new_n260_) & ((new_n242_ & ~new_n260_) | (~new_n242_ & new_n260_) | (~new_n243_ & (~new_n259_ | ((new_n262_ | (new_n241_ & ~new_n201_) | (~new_n241_ & new_n201_)) & (new_n245_ | (~new_n262_ & (~new_n241_ | new_n201_) & (new_n241_ | ~new_n201_)) | (new_n262_ & (~new_n241_ ^ ~new_n201_)))))));
  assign new_n241_ = new_n200_ ^ ~new_n208_;
  assign new_n242_ = (new_n196_ ^ ~new_n197_) ^ ((new_n198_ & ~new_n199_) | ((new_n198_ | ~new_n199_) & (~new_n198_ | new_n199_) & ((~new_n200_ & new_n208_) | (~new_n201_ & (new_n200_ | ~new_n208_) & (~new_n200_ | new_n208_)))));
  assign new_n243_ = ~new_n244_ & ((new_n198_ & ~new_n199_) | (~new_n198_ & new_n199_) | ((new_n200_ | ~new_n208_) & (new_n201_ | (~new_n200_ & new_n208_) | (new_n200_ & ~new_n208_)))) & ((new_n198_ ^ ~new_n199_) | (~new_n200_ & new_n208_) | (~new_n201_ & (new_n200_ | ~new_n208_) & (~new_n200_ | new_n208_)));
  assign new_n244_ = \a[14]  ^ (((\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[9]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[7]  | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n245_ = (new_n246_ | ~new_n247_) & ((new_n246_ & ~new_n247_) | (~new_n246_ & new_n247_) | ((~new_n248_ | new_n249_) & ((~new_n248_ & new_n249_) | (new_n248_ & ~new_n249_) | ((new_n250_ | ~new_n258_) & (new_n251_ | (~new_n250_ & new_n258_) | (new_n250_ & ~new_n258_))))));
  assign new_n246_ = \a[14]  ^ ((~new_n75_ | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[6]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[7]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[5]  | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n247_ = (new_n205_ | (~new_n206_ & new_n207_)) ^ (new_n204_ ^ (~\a[17]  ^ (new_n203_ & (~new_n66_ | ~new_n202_))));
  assign new_n248_ = new_n206_ ^ ~new_n207_;
  assign new_n249_ = \a[14]  ^ ((~new_n60_ | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[5]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[6]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[4]  | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n250_ = \a[14]  ^ ((~new_n63_ | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[4]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[5]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[3]  | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n251_ = (~new_n254_ | (\a[14]  ^ (new_n253_ & (~new_n66_ | ~new_n252_)))) & ((~new_n255_ & (new_n256_ | ~new_n257_)) | (new_n254_ & (~\a[14]  ^ (new_n253_ & (~new_n66_ | ~new_n252_)))) | (~new_n254_ & (~\a[14]  | ~new_n253_ | (new_n66_ & new_n252_)) & (\a[14]  | (new_n253_ & (~new_n66_ | ~new_n252_)))));
  assign new_n252_ = (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ) & (\a[13]  | \a[14] ) & (~\a[13]  | ~\a[14] );
  assign new_n253_ = (~\b[3]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[4]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & (~\b[2]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ));
  assign new_n254_ = ((\b[0]  & (\a[14]  ^ ~\a[15] ) & (\a[15]  | \a[16] ) & (~\a[15]  | ~\a[16] )) | (\b[1]  & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ) & (\a[16]  ^ ~\a[17] )) | ((\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ) & (\a[16]  | \a[17] ) & (~\a[16]  | ~\a[17] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[17]  & \b[0]  & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ));
  assign new_n255_ = \b[0]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] ) & (~\b[0]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[1]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & (~\b[1]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[0]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ));
  assign new_n256_ = \a[14]  ^ (((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & (~\b[2]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[1]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] )));
  assign new_n257_ = (\b[0]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) ^ ((~\b[0]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[1]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & (~\b[1]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[0]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] )));
  assign new_n258_ = (~\a[17]  | ((~\b[0]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[1]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[17]  & (~\b[0]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )))) ^ ((~\b[1]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[2]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  ^ ~\a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] )));
  assign new_n259_ = ~new_n244_ ^ ((new_n198_ ^ ~new_n199_) ^ ((~new_n200_ & new_n208_) | (~new_n201_ & (new_n200_ | ~new_n208_) & (~new_n200_ | new_n208_))));
  assign new_n260_ = \a[14]  ^ (new_n261_ & (~new_n252_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n261_ = (~\b[9]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[10]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & (~\b[8]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ));
  assign new_n262_ = \a[14]  ^ (((~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n80_ & (~\b[7]  ^ \b[8] )) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[7]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[8]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[6]  | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n263_ = ~new_n239_ ^ (new_n195_ ^ ~new_n238_);
  assign new_n264_ = ~new_n236_ ^ (new_n209_ ^ ((~new_n212_ & (new_n135_ | (~new_n134_ & new_n142_) | (new_n134_ & ~new_n142_)) & (~new_n135_ | (~new_n134_ ^ new_n142_))) | (~new_n195_ & (new_n212_ | (~new_n135_ & (new_n134_ | ~new_n142_) & (~new_n134_ | new_n142_)) | (new_n135_ & (new_n134_ ^ new_n142_))) & (~new_n212_ | (~new_n135_ ^ (~new_n134_ ^ new_n142_))))));
  assign new_n265_ = \a[14]  ^ ((~new_n149_ | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[12]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[13]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[11]  | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n266_ = new_n231_ & (~new_n214_ ^ (new_n187_ | (~new_n190_ & new_n213_)));
  assign new_n267_ = \a[14]  ^ (~\b[14]  | ((new_n164_ | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] ))));
  assign new_n268_ = \a[14]  ^ (((~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n114_ & (~\b[13]  ^ \b[14] )) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[13]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[14]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[12]  | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n269_ = ((\a[14]  & ((new_n54_ & \a[17] ) | (~new_n54_ & ~\a[17] ) | (~new_n176_ & (new_n177_ | ~new_n220_))) & ((new_n54_ ^ \a[17] ) | new_n176_ | (~new_n177_ & new_n220_))) | (~new_n270_ & (~\a[14]  | ((~new_n54_ | ~\a[17] ) & (new_n54_ | \a[17] ) & (new_n176_ | (~new_n177_ & new_n220_))) | ((~new_n54_ ^ \a[17] ) & ~new_n176_ & (new_n177_ | ~new_n220_))) & (\a[14]  | ((new_n54_ ^ \a[17] ) ^ (new_n176_ | (~new_n177_ & new_n220_)))))) ^ (\a[14]  ^ ((new_n174_ ^ \a[17] ) ^ ((new_n54_ & \a[17] ) | ((~new_n54_ | ~\a[17] ) & (new_n54_ | \a[17] ) & (new_n176_ | (~new_n177_ & new_n220_))))));
  assign new_n270_ = (~\a[14]  | (new_n177_ & ~new_n220_) | (~new_n177_ & new_n220_)) & (((~new_n223_ | ~\a[14] ) & ((new_n223_ & \a[14] ) | (~new_n223_ & ~\a[14] ) | ((~new_n225_ | ~\a[14] ) & (((~new_n226_ | ~\a[14] ) & (new_n228_ | (~new_n226_ & ~\a[14] ) | (new_n226_ & \a[14] ))) | (new_n225_ & \a[14] ) | (~new_n225_ & ~\a[14] ))))) | (\a[14]  & (~new_n177_ | new_n220_) & (new_n177_ | ~new_n220_)) | (~\a[14]  & (~new_n177_ ^ ~new_n220_)));
  assign new_n271_ = (~new_n272_ | ~\a[11] ) & ((~new_n272_ & ~\a[11] ) | (new_n272_ & \a[11] ) | ((~\a[11]  | ((~new_n223_ | ~\a[14] ) & (new_n223_ | \a[14] ) & ((new_n225_ & \a[14] ) | ((~new_n225_ | ~\a[14] ) & (new_n225_ | \a[14] ) & ((new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] )))))) | ((~new_n223_ ^ \a[14] ) & (~new_n225_ | ~\a[14] ) & ((new_n225_ & \a[14] ) | (~new_n225_ & ~\a[14] ) | ((~new_n226_ | ~\a[14] ) & (new_n228_ | (new_n226_ & \a[14] ) | (~new_n226_ & ~\a[14] )))))) & ((\a[11]  & ((new_n223_ & \a[14] ) | (~new_n223_ & ~\a[14] ) | ((~new_n225_ | ~\a[14] ) & ((new_n225_ & \a[14] ) | (~new_n225_ & ~\a[14] ) | ((~new_n226_ | ~\a[14] ) & (new_n228_ | (new_n226_ & \a[14] ) | (~new_n226_ & ~\a[14] )))))) & ((new_n223_ ^ \a[14] ) | (new_n225_ & \a[14] ) | ((~new_n225_ | ~\a[14] ) & (new_n225_ | \a[14] ) & ((new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] )))))) | (~\a[11]  & ((~new_n223_ ^ \a[14] ) ^ ((new_n225_ & \a[14] ) | ((~new_n225_ | ~\a[14] ) & (new_n225_ | \a[14] ) & ((new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] ))))))) | ((~\a[11]  | ((~new_n225_ | ~\a[14] ) & (new_n225_ | \a[14] ) & ((new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] )))) | ((~new_n225_ ^ \a[14] ) & (~new_n226_ | ~\a[14] ) & (new_n228_ | (new_n226_ & \a[14] ) | (~new_n226_ & ~\a[14] )))) & (new_n273_ | (\a[11]  & ((new_n225_ & \a[14] ) | (~new_n225_ & ~\a[14] ) | ((~new_n226_ | ~\a[14] ) & (new_n228_ | (new_n226_ & \a[14] ) | (~new_n226_ & ~\a[14] )))) & ((new_n225_ ^ \a[14] ) | (new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] )))) | (~\a[11]  & ((~new_n225_ ^ \a[14] ) ^ ((new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] ))))))))));
  assign new_n272_ = ((new_n223_ & \a[14] ) | ((~new_n223_ | ~\a[14] ) & (new_n223_ | \a[14] ) & ((new_n225_ & \a[14] ) | (((new_n226_ & \a[14] ) | (~new_n228_ & (new_n226_ | \a[14] ) & (~new_n226_ | ~\a[14] ))) & (~new_n225_ | ~\a[14] ) & (new_n225_ | \a[14] ))))) ^ (\a[14]  ^ (new_n177_ ^ ~new_n220_));
  assign new_n273_ = (~\a[11]  | (new_n275_ & ((new_n229_ & ~new_n267_) | (~new_n274_ & (new_n229_ | ~new_n267_) & (~new_n229_ | new_n267_)))) | (~new_n275_ & (~new_n229_ | new_n267_) & (new_n274_ | (~new_n229_ & new_n267_) | (new_n229_ & ~new_n267_)))) & (((~\a[11]  | (~new_n274_ & (new_n229_ | ~new_n267_) & (~new_n229_ | new_n267_)) | (new_n274_ & (new_n229_ ^ new_n267_))) & (((~new_n276_ | ~\a[11] ) & ((new_n276_ & \a[11] ) | (~new_n276_ & ~\a[11] ) | ((~new_n277_ | ~\a[11] ) & (new_n279_ | (new_n277_ & \a[11] ) | (~new_n277_ & ~\a[11] ))))) | (\a[11]  & (new_n274_ | (~new_n229_ & new_n267_) | (new_n229_ & ~new_n267_)) & (~new_n274_ | (~new_n229_ ^ new_n267_))) | (~\a[11]  & (new_n274_ ^ (~new_n229_ ^ new_n267_))))) | (\a[11]  & (~new_n275_ | ((~new_n229_ | new_n267_) & (new_n274_ | (~new_n229_ & new_n267_) | (new_n229_ & ~new_n267_)))) & (new_n275_ | (new_n229_ & ~new_n267_) | (~new_n274_ & (new_n229_ | ~new_n267_) & (~new_n229_ | new_n267_)))) | (~\a[11]  & (~new_n275_ ^ ((new_n229_ & ~new_n267_) | (~new_n274_ & (new_n229_ | ~new_n267_) & (~new_n229_ | new_n267_))))));
  assign new_n274_ = ~new_n230_ & (new_n230_ | new_n266_ | ((new_n268_ | (new_n190_ & ~new_n213_) | (~new_n190_ & new_n213_)) & (new_n232_ | (new_n268_ & (~new_n190_ ^ ~new_n213_)) | (~new_n268_ & (~new_n190_ | new_n213_) & (new_n190_ | ~new_n213_)))));
  assign new_n275_ = \a[14]  ^ (new_n182_ ^ ~new_n227_);
  assign new_n276_ = (~new_n230_ & ~new_n266_) ^ ((~new_n268_ & (~new_n190_ | new_n213_) & (new_n190_ | ~new_n213_)) | (~new_n232_ & (~new_n268_ | (new_n190_ ^ ~new_n213_)) & (new_n268_ | (new_n190_ & ~new_n213_) | (~new_n190_ & new_n213_))));
  assign new_n277_ = new_n232_ ^ ~new_n278_;
  assign new_n278_ = ~new_n268_ ^ (new_n190_ ^ ~new_n213_);
  assign new_n279_ = (~new_n280_ | new_n318_) & ((new_n280_ & ~new_n318_) | (~new_n280_ & new_n318_) | (~new_n281_ & (((new_n319_ | (~new_n240_ & new_n263_) | (new_n240_ & ~new_n263_)) & (new_n283_ | (~new_n319_ & (new_n240_ | ~new_n263_) & (~new_n240_ | new_n263_)) | (new_n319_ & (new_n240_ ^ new_n263_)))) | new_n281_ | new_n317_)));
  assign new_n280_ = (new_n235_ | (new_n264_ & (new_n237_ | (~new_n240_ & new_n263_)))) ^ (new_n233_ ^ ~new_n265_);
  assign new_n281_ = ~new_n282_ & (~new_n264_ | (~new_n237_ & (new_n240_ | ~new_n263_))) & (new_n264_ | new_n237_ | (~new_n240_ & new_n263_));
  assign new_n282_ = \a[11]  ^ (((\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\b[14]  ^ ((\b[13]  & \b[14] ) | (~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] ))))) & (~\b[14]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[13]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n283_ = (~new_n284_ | new_n316_) & ((~new_n286_ & (~new_n315_ | (~new_n288_ & (new_n291_ | ~new_n314_)))) | (new_n284_ & ~new_n316_) | (~new_n284_ & new_n316_));
  assign new_n284_ = new_n285_ ^ (new_n243_ | (new_n259_ & ((~new_n262_ & (new_n201_ | (~new_n200_ & new_n208_) | (new_n200_ & ~new_n208_)) & (~new_n201_ | (~new_n200_ ^ new_n208_))) | (~new_n245_ & (new_n262_ | (~new_n201_ & (new_n200_ | ~new_n208_) & (~new_n200_ | new_n208_)) | (new_n201_ & (new_n200_ ^ new_n208_))) & (~new_n262_ | (~new_n201_ ^ (~new_n200_ ^ new_n208_)))))));
  assign new_n285_ = ~new_n260_ ^ ((new_n196_ ^ ~new_n197_) ^ ((new_n198_ & ~new_n199_) | ((new_n198_ | ~new_n199_) & (~new_n198_ | new_n199_) & ((~new_n200_ & new_n208_) | (~new_n201_ & (new_n200_ | ~new_n208_) & (~new_n200_ | new_n208_))))));
  assign new_n286_ = ~new_n287_ & (~new_n259_ | ((new_n262_ | (~new_n201_ & (new_n200_ | ~new_n208_) & (~new_n200_ | new_n208_)) | (new_n201_ & (new_n200_ ^ new_n208_))) & (new_n245_ | (~new_n262_ & (new_n201_ | (~new_n200_ & new_n208_) | (new_n200_ & ~new_n208_)) & (~new_n201_ | (~new_n200_ ^ new_n208_))) | (new_n262_ & (new_n201_ ^ (~new_n200_ ^ new_n208_)))))) & (new_n259_ | (~new_n262_ & (new_n201_ | (~new_n200_ & new_n208_) | (new_n200_ & ~new_n208_)) & (~new_n201_ | (~new_n200_ ^ new_n208_))) | (~new_n245_ & (new_n262_ | (~new_n201_ & (new_n200_ | ~new_n208_) & (~new_n200_ | new_n208_)) | (new_n201_ & (new_n200_ ^ new_n208_))) & (~new_n262_ | (~new_n201_ ^ (~new_n200_ ^ new_n208_)))));
  assign new_n287_ = \a[11]  ^ ((~new_n106_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[11]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[12]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[10]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n288_ = ~new_n290_ & (~new_n245_ | new_n289_) & (new_n245_ | ~new_n289_);
  assign new_n289_ = ~new_n262_ ^ (~new_n201_ ^ (new_n200_ ^ ~new_n208_));
  assign new_n290_ = \a[11]  ^ ((~new_n112_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[10]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[11]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[9]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n291_ = (~new_n293_ | new_n311_) & ((new_n293_ & ~new_n311_) | (~new_n293_ & new_n311_) | (~new_n294_ & (~new_n310_ | ((new_n313_ | (new_n292_ & ~new_n251_) | (~new_n292_ & new_n251_)) & (new_n296_ | (~new_n313_ & (~new_n292_ | new_n251_) & (new_n292_ | ~new_n251_)) | (new_n313_ & (~new_n292_ ^ ~new_n251_)))))));
  assign new_n292_ = new_n250_ ^ ~new_n258_;
  assign new_n293_ = (new_n246_ ^ ~new_n247_) ^ ((new_n248_ & ~new_n249_) | ((new_n248_ | ~new_n249_) & (~new_n248_ | new_n249_) & ((~new_n250_ & new_n258_) | (~new_n251_ & (new_n250_ | ~new_n258_) & (~new_n250_ | new_n258_)))));
  assign new_n294_ = ~new_n295_ & ((new_n248_ & ~new_n249_) | (~new_n248_ & new_n249_) | ((new_n250_ | ~new_n258_) & (new_n251_ | (~new_n250_ & new_n258_) | (new_n250_ & ~new_n258_)))) & ((new_n248_ ^ ~new_n249_) | (~new_n250_ & new_n258_) | (~new_n251_ & (new_n250_ | ~new_n258_) & (~new_n250_ | new_n258_)));
  assign new_n295_ = \a[11]  ^ (((\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[9]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[7]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n296_ = (new_n297_ | ~new_n298_) & ((new_n297_ & ~new_n298_) | (~new_n297_ & new_n298_) | ((~new_n299_ | new_n300_) & ((~new_n299_ & new_n300_) | (new_n299_ & ~new_n300_) | ((new_n301_ | ~new_n309_) & (new_n302_ | (~new_n301_ & new_n309_) | (new_n301_ & ~new_n309_))))));
  assign new_n297_ = \a[11]  ^ ((~new_n75_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[6]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[7]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[5]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n298_ = (new_n255_ | (~new_n256_ & new_n257_)) ^ (new_n254_ ^ (~\a[14]  ^ (new_n253_ & (~new_n66_ | ~new_n252_))));
  assign new_n299_ = new_n256_ ^ ~new_n257_;
  assign new_n300_ = \a[11]  ^ ((~new_n60_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[5]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[6]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[4]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n301_ = \a[11]  ^ ((~new_n63_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[4]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[5]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[3]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n302_ = (~new_n305_ | (\a[11]  ^ (new_n304_ & (~new_n66_ | ~new_n303_)))) & ((~new_n306_ & (new_n307_ | ~new_n308_)) | (new_n305_ & (~\a[11]  ^ (new_n304_ & (~new_n66_ | ~new_n303_)))) | (~new_n305_ & (~\a[11]  | ~new_n304_ | (new_n66_ & new_n303_)) & (\a[11]  | (new_n304_ & (~new_n66_ | ~new_n303_)))));
  assign new_n303_ = (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] );
  assign new_n304_ = (~\b[3]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[4]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[2]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ));
  assign new_n305_ = ((\b[0]  & (\a[11]  ^ ~\a[12] ) & (\a[12]  | \a[13] ) & (~\a[12]  | ~\a[13] )) | (\b[1]  & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ) & (\a[13]  ^ ~\a[14] )) | ((\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ) & (\a[13]  | \a[14] ) & (~\a[13]  | ~\a[14] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[14]  & \b[0]  & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ));
  assign new_n306_ = \b[0]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] ) & (~\b[0]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[1]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[0]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ));
  assign new_n307_ = \a[11]  ^ (((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[2]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] )));
  assign new_n308_ = (\b[0]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] )) ^ ((~\b[0]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[1]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[0]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] )));
  assign new_n309_ = (~\a[14]  | ((~\b[0]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[1]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )))) ^ ((~\b[1]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[2]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  ^ ~\a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[12]  ^ ~\a[13] ) | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] )));
  assign new_n310_ = ~new_n295_ ^ ((new_n248_ ^ ~new_n249_) ^ ((~new_n250_ & new_n258_) | (~new_n251_ & (new_n250_ | ~new_n258_) & (~new_n250_ | new_n258_))));
  assign new_n311_ = \a[11]  ^ (new_n312_ & (~new_n303_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n312_ = (~\b[9]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[10]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[8]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ));
  assign new_n313_ = \a[11]  ^ (((~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n80_ & (~\b[7]  ^ \b[8] )) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[7]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[8]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[6]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n314_ = ~new_n290_ ^ (new_n245_ ^ ~new_n289_);
  assign new_n315_ = ~new_n287_ ^ (new_n259_ ^ ((~new_n262_ & (new_n201_ | (~new_n200_ & new_n208_) | (new_n200_ & ~new_n208_)) & (~new_n201_ | (~new_n200_ ^ new_n208_))) | (~new_n245_ & (new_n262_ | (~new_n201_ & (new_n200_ | ~new_n208_) & (~new_n200_ | new_n208_)) | (new_n201_ & (new_n200_ ^ new_n208_))) & (~new_n262_ | (~new_n201_ ^ (~new_n200_ ^ new_n208_))))));
  assign new_n316_ = \a[11]  ^ ((~new_n149_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[12]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[13]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[11]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n317_ = new_n282_ & (~new_n264_ ^ (new_n237_ | (~new_n240_ & new_n263_)));
  assign new_n318_ = \a[11]  ^ (~\b[14]  | ((new_n164_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] ))));
  assign new_n319_ = \a[11]  ^ (((~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n114_ & (~\b[13]  ^ \b[14] )) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[13]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[14]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[12]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n320_ = \a[14]  ^ ((new_n176_ | (~new_n177_ & new_n220_)) ^ (new_n54_ ^ \a[17] ));
  assign new_n321_ = \a[8]  & ((new_n269_ & \a[11] ) | (~new_n269_ & ~\a[11] ) | ((~\a[11]  | (~new_n270_ & new_n320_) | (new_n270_ & ~new_n320_)) & (new_n271_ | (\a[11]  & (new_n270_ | ~new_n320_) & (~new_n270_ | new_n320_)) | (~\a[11]  & (new_n270_ ^ new_n320_))))) & ((new_n269_ ^ \a[11] ) | (\a[11]  & (new_n270_ | ~new_n320_) & (~new_n270_ | new_n320_)) | (~new_n271_ & (~\a[11]  | (~new_n270_ & new_n320_) | (new_n270_ & ~new_n320_)) & (\a[11]  | (~new_n270_ ^ new_n320_))));
  assign new_n322_ = (~\a[8]  | (new_n271_ & ~new_n323_) | (~new_n271_ & new_n323_)) & (((~new_n324_ | ~\a[8] ) & ((new_n324_ & \a[8] ) | (~new_n324_ & ~\a[8] ) | ((~new_n325_ | ~\a[8] ) & (((~new_n326_ | ~\a[8] ) & (new_n328_ | (~new_n326_ & ~\a[8] ) | (new_n326_ & \a[8] ))) | (new_n325_ & \a[8] ) | (~new_n325_ & ~\a[8] ))))) | (\a[8]  & (~new_n271_ | new_n323_) & (new_n271_ | ~new_n323_)) | (~\a[8]  & (~new_n271_ ^ ~new_n323_)));
  assign new_n323_ = \a[11]  ^ (new_n270_ ^ ~new_n320_);
  assign new_n324_ = (~new_n272_ ^ ~\a[11] ) ^ ((\a[11]  & ((new_n223_ & \a[14] ) | (~new_n223_ & ~\a[14] ) | ((~new_n225_ | ~\a[14] ) & ((new_n225_ & \a[14] ) | (~new_n225_ & ~\a[14] ) | ((~new_n226_ | ~\a[14] ) & (new_n228_ | (new_n226_ & \a[14] ) | (~new_n226_ & ~\a[14] )))))) & ((new_n223_ ^ \a[14] ) | (new_n225_ & \a[14] ) | ((~new_n225_ | ~\a[14] ) & (new_n225_ | \a[14] ) & ((new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] )))))) | ((~\a[11]  | ((~new_n223_ | ~\a[14] ) & (new_n223_ | \a[14] ) & ((new_n225_ & \a[14] ) | ((~new_n225_ | ~\a[14] ) & (new_n225_ | \a[14] ) & ((new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] )))))) | ((~new_n223_ ^ \a[14] ) & (~new_n225_ | ~\a[14] ) & ((new_n225_ & \a[14] ) | (~new_n225_ & ~\a[14] ) | ((~new_n226_ | ~\a[14] ) & (new_n228_ | (new_n226_ & \a[14] ) | (~new_n226_ & ~\a[14] )))))) & (\a[11]  | ((new_n223_ ^ \a[14] ) ^ ((new_n225_ & \a[14] ) | ((~new_n225_ | ~\a[14] ) & (new_n225_ | \a[14] ) & ((new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] ))))))) & ((\a[11]  & ((new_n225_ & \a[14] ) | (~new_n225_ & ~\a[14] ) | ((~new_n226_ | ~\a[14] ) & (new_n228_ | (new_n226_ & \a[14] ) | (~new_n226_ & ~\a[14] )))) & ((new_n225_ ^ \a[14] ) | (new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] )))) | (~new_n273_ & (~\a[11]  | ((~new_n225_ | ~\a[14] ) & (new_n225_ | \a[14] ) & ((new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] )))) | ((~new_n225_ ^ \a[14] ) & (~new_n226_ | ~\a[14] ) & (new_n228_ | (new_n226_ & \a[14] ) | (~new_n226_ & ~\a[14] )))) & (\a[11]  | ((new_n225_ ^ \a[14] ) ^ ((new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] )))))))));
  assign new_n325_ = ((\a[11]  & ((new_n225_ & \a[14] ) | (~new_n225_ & ~\a[14] ) | ((~new_n226_ | ~\a[14] ) & (new_n228_ | (new_n226_ & \a[14] ) | (~new_n226_ & ~\a[14] )))) & ((new_n225_ ^ \a[14] ) | (new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] )))) | (~new_n273_ & (~\a[11]  | ((~new_n225_ | ~\a[14] ) & (new_n225_ | \a[14] ) & ((new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] )))) | ((~new_n225_ ^ \a[14] ) & (~new_n226_ | ~\a[14] ) & (new_n228_ | (new_n226_ & \a[14] ) | (~new_n226_ & ~\a[14] )))) & (\a[11]  | ((new_n225_ ^ \a[14] ) ^ ((new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] ))))))) ^ (\a[11]  ^ (((new_n225_ & \a[14] ) | ((~new_n225_ | ~\a[14] ) & (new_n225_ | \a[14] ) & ((new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] ))))) ^ (new_n223_ ^ \a[14] )));
  assign new_n326_ = new_n273_ ^ ~new_n327_;
  assign new_n327_ = \a[11]  ^ ((new_n225_ ^ \a[14] ) ^ ((new_n226_ & \a[14] ) | (~new_n228_ & (~new_n226_ | ~\a[14] ) & (new_n226_ | \a[14] ))));
  assign new_n328_ = (~new_n330_ | ~\a[8] ) & ((new_n330_ & \a[8] ) | (~new_n330_ & ~\a[8] ) | ((~\a[8]  | (((new_n276_ & \a[11] ) | ((~new_n276_ | ~\a[11] ) & (new_n276_ | \a[11] ) & ((new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] ))))) & (~new_n329_ | ~\a[11] ) & (new_n329_ | \a[11] )) | ((~new_n276_ | ~\a[11] ) & ((new_n276_ & \a[11] ) | (~new_n276_ & ~\a[11] ) | ((~new_n277_ | ~\a[11] ) & (new_n279_ | (new_n277_ & \a[11] ) | (~new_n277_ & ~\a[11] )))) & (~new_n329_ ^ \a[11] ))) & ((\a[8]  & (((~new_n276_ | ~\a[11] ) & ((new_n276_ & \a[11] ) | (~new_n276_ & ~\a[11] ) | ((~new_n277_ | ~\a[11] ) & (new_n279_ | (new_n277_ & \a[11] ) | (~new_n277_ & ~\a[11] ))))) | (new_n329_ & \a[11] ) | (~new_n329_ & ~\a[11] )) & ((new_n276_ & \a[11] ) | ((~new_n276_ | ~\a[11] ) & (new_n276_ | \a[11] ) & ((new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] )))) | (new_n329_ ^ \a[11] ))) | (~\a[8]  & (((~new_n276_ | ~\a[11] ) & ((new_n276_ & \a[11] ) | (~new_n276_ & ~\a[11] ) | ((~new_n277_ | ~\a[11] ) & (new_n279_ | (new_n277_ & \a[11] ) | (~new_n277_ & ~\a[11] ))))) ^ (new_n329_ ^ \a[11] ))) | ((~\a[8]  | ((~new_n276_ | ~\a[11] ) & (new_n276_ | \a[11] ) & ((new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] )))) | ((~new_n276_ ^ \a[11] ) & (~new_n277_ | ~\a[11] ) & (new_n279_ | (new_n277_ & \a[11] ) | (~new_n277_ & ~\a[11] )))) & (new_n331_ | (\a[8]  & ((new_n276_ & \a[11] ) | (~new_n276_ & ~\a[11] ) | ((~new_n277_ | ~\a[11] ) & (new_n279_ | (new_n277_ & \a[11] ) | (~new_n277_ & ~\a[11] )))) & ((new_n276_ ^ \a[11] ) | (new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] )))) | (~\a[8]  & ((~new_n276_ ^ \a[11] ) ^ ((new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] ))))))))));
  assign new_n329_ = ~new_n274_ ^ (~new_n229_ ^ new_n267_);
  assign new_n330_ = ((\a[11]  & (new_n274_ | (~new_n229_ & new_n267_) | (new_n229_ & ~new_n267_)) & (~new_n274_ | (~new_n229_ ^ new_n267_))) | (((new_n276_ & \a[11] ) | ((~new_n276_ | ~\a[11] ) & (new_n276_ | \a[11] ) & ((new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] ))))) & (~\a[11]  | (~new_n274_ & (new_n229_ | ~new_n267_) & (~new_n229_ | new_n267_)) | (new_n274_ & (new_n229_ ^ new_n267_))) & (\a[11]  | (~new_n274_ ^ (~new_n229_ ^ new_n267_))))) ^ (\a[11]  ^ (new_n275_ ^ ((new_n229_ & ~new_n267_) | (~new_n274_ & (new_n229_ | ~new_n267_) & (~new_n229_ | new_n267_)))));
  assign new_n331_ = (~\a[8]  | (new_n333_ & ((new_n280_ & ~new_n318_) | (~new_n332_ & (new_n280_ | ~new_n318_) & (~new_n280_ | new_n318_)))) | (~new_n333_ & (~new_n280_ | new_n318_) & (new_n332_ | (~new_n280_ & new_n318_) | (new_n280_ & ~new_n318_)))) & (((~\a[8]  | (~new_n332_ & (new_n280_ | ~new_n318_) & (~new_n280_ | new_n318_)) | (new_n332_ & (new_n280_ ^ new_n318_))) & (((~new_n334_ | ~\a[8] ) & ((new_n334_ & \a[8] ) | (~new_n334_ & ~\a[8] ) | ((~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] ))))) | (\a[8]  & (new_n332_ | (~new_n280_ & new_n318_) | (new_n280_ & ~new_n318_)) & (~new_n332_ | (~new_n280_ ^ new_n318_))) | (~\a[8]  & (new_n332_ ^ (~new_n280_ ^ new_n318_))))) | (\a[8]  & (~new_n333_ | ((~new_n280_ | new_n318_) & (new_n332_ | (~new_n280_ & new_n318_) | (new_n280_ & ~new_n318_)))) & (new_n333_ | (new_n280_ & ~new_n318_) | (~new_n332_ & (new_n280_ | ~new_n318_) & (~new_n280_ | new_n318_)))) | (~\a[8]  & (~new_n333_ ^ ((new_n280_ & ~new_n318_) | (~new_n332_ & (new_n280_ | ~new_n318_) & (~new_n280_ | new_n318_))))));
  assign new_n332_ = ~new_n281_ & (new_n281_ | new_n317_ | ((new_n319_ | (new_n240_ & ~new_n263_) | (~new_n240_ & new_n263_)) & (new_n283_ | (new_n319_ & (~new_n240_ ^ ~new_n263_)) | (~new_n319_ & (~new_n240_ | new_n263_) & (new_n240_ | ~new_n263_)))));
  assign new_n333_ = \a[11]  ^ (new_n232_ ^ ~new_n278_);
  assign new_n334_ = (~new_n281_ & ~new_n317_) ^ ((~new_n319_ & (~new_n240_ | new_n263_) & (new_n240_ | ~new_n263_)) | (~new_n283_ & (~new_n319_ | (new_n240_ ^ ~new_n263_)) & (new_n319_ | (new_n240_ & ~new_n263_) | (~new_n240_ & new_n263_))));
  assign new_n335_ = new_n283_ ^ ~new_n336_;
  assign new_n336_ = ~new_n319_ ^ (new_n240_ ^ ~new_n263_);
  assign new_n337_ = (~new_n338_ | new_n376_) & ((new_n338_ & ~new_n376_) | (~new_n338_ & new_n376_) | (~new_n339_ & (((new_n377_ | (~new_n291_ & new_n314_) | (new_n291_ & ~new_n314_)) & (new_n341_ | (~new_n377_ & (new_n291_ | ~new_n314_) & (~new_n291_ | new_n314_)) | (new_n377_ & (new_n291_ ^ new_n314_)))) | new_n339_ | new_n375_)));
  assign new_n338_ = (new_n286_ | (new_n315_ & (new_n288_ | (~new_n291_ & new_n314_)))) ^ (new_n284_ ^ ~new_n316_);
  assign new_n339_ = ~new_n340_ & (~new_n315_ | (~new_n288_ & (new_n291_ | ~new_n314_))) & (new_n315_ | new_n288_ | (~new_n291_ & new_n314_));
  assign new_n340_ = \a[8]  ^ (((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\b[14]  ^ ((\b[13]  & \b[14] ) | (~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] ))))) & (~\b[14]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[13]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n341_ = (~new_n342_ | new_n374_) & ((~new_n344_ & (~new_n373_ | (~new_n346_ & (new_n349_ | ~new_n372_)))) | (new_n342_ & ~new_n374_) | (~new_n342_ & new_n374_));
  assign new_n342_ = new_n343_ ^ (new_n294_ | (new_n310_ & ((~new_n313_ & (new_n251_ | (~new_n250_ & new_n258_) | (new_n250_ & ~new_n258_)) & (~new_n251_ | (~new_n250_ ^ new_n258_))) | (~new_n296_ & (new_n313_ | (~new_n251_ & (new_n250_ | ~new_n258_) & (~new_n250_ | new_n258_)) | (new_n251_ & (new_n250_ ^ new_n258_))) & (~new_n313_ | (~new_n251_ ^ (~new_n250_ ^ new_n258_)))))));
  assign new_n343_ = ~new_n311_ ^ ((new_n246_ ^ ~new_n247_) ^ ((new_n248_ & ~new_n249_) | ((new_n248_ | ~new_n249_) & (~new_n248_ | new_n249_) & ((~new_n250_ & new_n258_) | (~new_n251_ & (new_n250_ | ~new_n258_) & (~new_n250_ | new_n258_))))));
  assign new_n344_ = ~new_n345_ & (~new_n310_ | ((new_n313_ | (~new_n251_ & (new_n250_ | ~new_n258_) & (~new_n250_ | new_n258_)) | (new_n251_ & (new_n250_ ^ new_n258_))) & (new_n296_ | (~new_n313_ & (new_n251_ | (~new_n250_ & new_n258_) | (new_n250_ & ~new_n258_)) & (~new_n251_ | (~new_n250_ ^ new_n258_))) | (new_n313_ & (new_n251_ ^ (~new_n250_ ^ new_n258_)))))) & (new_n310_ | (~new_n313_ & (new_n251_ | (~new_n250_ & new_n258_) | (new_n250_ & ~new_n258_)) & (~new_n251_ | (~new_n250_ ^ new_n258_))) | (~new_n296_ & (new_n313_ | (~new_n251_ & (new_n250_ | ~new_n258_) & (~new_n250_ | new_n258_)) | (new_n251_ & (new_n250_ ^ new_n258_))) & (~new_n313_ | (~new_n251_ ^ (~new_n250_ ^ new_n258_)))));
  assign new_n345_ = \a[8]  ^ ((~new_n106_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[11]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[12]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[10]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n346_ = ~new_n348_ & (~new_n296_ | new_n347_) & (new_n296_ | ~new_n347_);
  assign new_n347_ = ~new_n313_ ^ (~new_n251_ ^ (new_n250_ ^ ~new_n258_));
  assign new_n348_ = \a[8]  ^ ((~new_n112_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[10]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[11]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[9]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n349_ = (~new_n351_ | new_n369_) & ((new_n351_ & ~new_n369_) | (~new_n351_ & new_n369_) | (~new_n352_ & (~new_n368_ | ((new_n371_ | (new_n350_ & ~new_n302_) | (~new_n350_ & new_n302_)) & (new_n354_ | (~new_n371_ & (~new_n350_ | new_n302_) & (new_n350_ | ~new_n302_)) | (new_n371_ & (~new_n350_ ^ ~new_n302_)))))));
  assign new_n350_ = new_n301_ ^ ~new_n309_;
  assign new_n351_ = (new_n297_ ^ ~new_n298_) ^ ((new_n299_ & ~new_n300_) | ((new_n299_ | ~new_n300_) & (~new_n299_ | new_n300_) & ((~new_n301_ & new_n309_) | (~new_n302_ & (new_n301_ | ~new_n309_) & (~new_n301_ | new_n309_)))));
  assign new_n352_ = ~new_n353_ & ((new_n299_ & ~new_n300_) | (~new_n299_ & new_n300_) | ((new_n301_ | ~new_n309_) & (new_n302_ | (~new_n301_ & new_n309_) | (new_n301_ & ~new_n309_)))) & ((new_n299_ ^ ~new_n300_) | (~new_n301_ & new_n309_) | (~new_n302_ & (new_n301_ | ~new_n309_) & (~new_n301_ | new_n309_)));
  assign new_n353_ = \a[8]  ^ (((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[9]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[7]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n354_ = (~new_n355_ | new_n356_) & ((new_n355_ & ~new_n356_) | (~new_n355_ & new_n356_) | ((~new_n357_ | new_n358_) & ((~new_n357_ & new_n358_) | (new_n357_ & ~new_n358_) | ((new_n359_ | ~new_n367_) & (new_n360_ | (~new_n359_ & new_n367_) | (new_n359_ & ~new_n367_))))));
  assign new_n355_ = (new_n306_ | (~new_n307_ & new_n308_)) ^ (new_n305_ ^ (~\a[11]  ^ (new_n304_ & (~new_n66_ | ~new_n303_))));
  assign new_n356_ = \a[8]  ^ ((~new_n75_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[6]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[7]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[5]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n357_ = new_n307_ ^ ~new_n308_;
  assign new_n358_ = \a[8]  ^ ((~new_n60_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[5]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[6]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[4]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n359_ = \a[8]  ^ ((~new_n63_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[4]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[5]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[3]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n360_ = (~new_n363_ | (\a[8]  ^ (new_n362_ & (~new_n66_ | ~new_n361_)))) & ((~new_n364_ & (new_n365_ | ~new_n366_)) | (new_n363_ & (~\a[8]  ^ (new_n362_ & (~new_n66_ | ~new_n361_)))) | (~new_n363_ & (~\a[8]  | ~new_n362_ | (new_n66_ & new_n361_)) & (\a[8]  | (new_n362_ & (~new_n66_ | ~new_n361_)))));
  assign new_n361_ = (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] );
  assign new_n362_ = (~\b[3]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[4]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[2]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ));
  assign new_n363_ = ((\b[0]  & (\a[8]  ^ ~\a[9] ) & (\a[9]  | \a[10] ) & (~\a[9]  | ~\a[10] )) | (\b[1]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  ^ ~\a[11] )) | ((\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[11]  & \b[0]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ));
  assign new_n364_ = \b[0]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] ) & (~\b[0]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[1]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ));
  assign new_n365_ = \a[8]  ^ (((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[2]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )));
  assign new_n366_ = (\b[0]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] )) ^ ((~\b[0]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[1]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )));
  assign new_n367_ = (~\a[11]  | ((~\b[0]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )))) ^ ((~\b[1]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[2]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[9]  ^ ~\a[10] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] )));
  assign new_n368_ = ~new_n353_ ^ ((new_n299_ ^ ~new_n300_) ^ ((~new_n301_ & new_n309_) | (~new_n302_ & (new_n301_ | ~new_n309_) & (~new_n301_ | new_n309_))));
  assign new_n369_ = \a[8]  ^ (new_n370_ & (~new_n361_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n370_ = (~\b[9]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[10]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[8]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ));
  assign new_n371_ = \a[8]  ^ (((~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n80_ & (~\b[7]  ^ \b[8] )) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[7]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[8]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[6]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n372_ = ~new_n348_ ^ (new_n296_ ^ ~new_n347_);
  assign new_n373_ = ~new_n345_ ^ (new_n310_ ^ ((~new_n313_ & (new_n251_ | (~new_n250_ & new_n258_) | (new_n250_ & ~new_n258_)) & (~new_n251_ | (~new_n250_ ^ new_n258_))) | (~new_n296_ & (new_n313_ | (~new_n251_ & (new_n250_ | ~new_n258_) & (~new_n250_ | new_n258_)) | (new_n251_ & (new_n250_ ^ new_n258_))) & (~new_n313_ | (~new_n251_ ^ (~new_n250_ ^ new_n258_))))));
  assign new_n374_ = \a[8]  ^ ((~new_n149_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[12]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[13]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[11]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n375_ = new_n340_ & (~new_n315_ ^ (new_n288_ | (~new_n291_ & new_n314_)));
  assign new_n376_ = \a[8]  ^ (~\b[14]  | ((new_n164_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] ))));
  assign new_n377_ = \a[8]  ^ (((~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n114_ & (~\b[13]  ^ \b[14] )) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[13]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[14]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[12]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n378_ = \a[8]  ^ ((new_n269_ ^ \a[11] ) ^ ((\a[11]  & (new_n270_ | ~new_n320_) & (~new_n270_ | new_n320_)) | (~new_n271_ & (~\a[11]  | (~new_n270_ & new_n320_) | (new_n270_ & ~new_n320_)) & (\a[11]  | (~new_n270_ ^ new_n320_)))));
  assign new_n379_ = (new_n413_ ^ \a[14] ) ^ ((new_n380_ & \a[14] ) | ((new_n380_ | \a[14] ) & (~new_n380_ | ~\a[14] ) & ((new_n409_ & \a[14] ) | ((new_n410_ | (~new_n411_ & new_n412_)) & (~new_n409_ | ~\a[14] ) & (new_n409_ | \a[14] )))));
  assign new_n380_ = (new_n381_ ^ \a[17] ) ^ ((new_n405_ & \a[17] ) | ((~new_n405_ | ~\a[17] ) & (new_n405_ | \a[17] ) & ((~new_n407_ & new_n408_) | (new_n406_ & \a[17] ))));
  assign new_n381_ = (~new_n382_ ^ \a[20] ) ^ ((~new_n403_ | ~\a[20] ) & ((new_n403_ & \a[20] ) | (~new_n403_ & ~\a[20] ) | ((~new_n404_ | ~\a[20] ) & (((~new_n166_ | ~\a[20] ) & (new_n154_ | (new_n166_ & \a[20] ) | (~new_n166_ & ~\a[20] ))) | (new_n404_ & \a[20] ) | (~new_n404_ & ~\a[20] )))));
  assign new_n382_ = ~new_n398_ ^ ((~new_n383_ | new_n402_) & ((new_n383_ & ~new_n402_) | (~new_n383_ & new_n402_) | (~new_n392_ & (~new_n397_ | (~new_n394_ & ~new_n396_)))));
  assign new_n383_ = new_n390_ ^ (new_n384_ | (new_n387_ & ~new_n388_));
  assign new_n384_ = ~new_n386_ & (new_n385_ ^ ~\a[26] );
  assign new_n385_ = (~\b[10]  | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (~\a[24]  ^ ~\a[25] ) | (~\a[23]  ^ ~\a[24] )) & (~\b[11]  | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] ) | (~\a[23]  ^ ~\a[24] )) & (~\b[12]  | (\a[25]  ^ \a[26] ) | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~new_n106_ | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ));
  assign new_n386_ = (~\b[8]  | ~\a[27]  | (\a[26]  & ~\a[27] ) | (~\a[26]  & \a[27] )) & (~\b[9]  | (\a[26]  ^ ~\a[27] ));
  assign new_n387_ = ~new_n386_ ^ (new_n385_ ^ ~\a[26] );
  assign new_n388_ = ~new_n389_ & (~new_n170_ | ((new_n169_ | new_n161_) & ((new_n169_ & new_n161_) | (~new_n169_ & ~new_n161_) | ((new_n107_ | new_n109_) & ((new_n107_ & new_n109_) | (~new_n107_ & ~new_n109_) | (~new_n100_ & ~new_n108_))))));
  assign new_n389_ = (new_n171_ ^ ~\a[26] ) & ((\b[8]  & (\a[26]  ^ \a[27] )) | (\b[7]  & \a[27]  & (\a[26]  | ~\a[27] ) & (~\a[26]  | \a[27] )));
  assign new_n390_ = (new_n391_ ^ ~\a[26] ) ^ ((\b[10]  & (\a[26]  ^ \a[27] )) | (\b[9]  & \a[27]  & (\a[26]  | ~\a[27] ) & (~\a[26]  | \a[27] )));
  assign new_n391_ = (~\b[11]  | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (~\a[24]  ^ ~\a[25] ) | (~\a[23]  ^ ~\a[24] )) & (~\b[12]  | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] ) | (~\a[23]  ^ ~\a[24] )) & (~\b[13]  | (\a[25]  ^ \a[26] ) | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~new_n149_ | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ));
  assign new_n392_ = ~new_n393_ & (~new_n387_ | new_n388_) & (new_n387_ | ~new_n388_);
  assign new_n393_ = \a[23]  ^ (((\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (~\b[14]  ^ ((\b[13]  & \b[14] ) | (~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] ))))) & (~\b[13]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[21]  ^ ~\a[22] ) | (~\a[20]  ^ ~\a[21] )) & (~\b[14]  | (~\a[21]  & ~\a[22] ) | (\a[21]  & \a[22] ) | (~\a[20]  ^ ~\a[21] )));
  assign new_n394_ = ~new_n173_ & (~new_n395_ | new_n170_) & (new_n395_ | ~new_n170_);
  assign new_n395_ = (new_n169_ | new_n161_) & (~new_n158_ | ((new_n107_ | new_n109_) & ((~new_n100_ & ~new_n108_) | (new_n107_ & new_n109_) | (~new_n107_ & ~new_n109_))));
  assign new_n396_ = new_n168_ & (new_n167_ | (new_n157_ & (new_n156_ | (new_n99_ & ((new_n110_ & ~new_n111_) | (~new_n56_ & (~new_n110_ | new_n111_) & (new_n110_ | ~new_n111_)))))));
  assign new_n397_ = ~new_n393_ ^ (new_n387_ ^ ~new_n388_);
  assign new_n398_ = \a[23]  ^ (new_n400_ ^ (new_n399_ | (new_n390_ & (new_n384_ | (new_n387_ & ~new_n388_)))));
  assign new_n399_ = (new_n391_ ^ ~\a[26] ) & ((\b[10]  & (\a[26]  ^ \a[27] )) | (\b[9]  & \a[27]  & (\a[26]  | ~\a[27] ) & (~\a[26]  | \a[27] )));
  assign new_n400_ = (new_n401_ ^ ~\a[26] ) ^ ((\b[11]  & (\a[26]  ^ \a[27] )) | (\b[10]  & \a[27]  & (\a[26]  | ~\a[27] ) & (~\a[26]  | \a[27] )));
  assign new_n401_ = ((~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n114_ & (~\b[13]  ^ \b[14] )) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~\b[12]  | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (~\a[24]  ^ ~\a[25] ) | (~\a[23]  ^ ~\a[24] )) & (~\b[13]  | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] ) | (~\a[23]  ^ ~\a[24] )) & (~\b[14]  | (\a[25]  ^ \a[26] ) | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ));
  assign new_n402_ = \a[23]  ^ (~\b[14]  | (((\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[21]  ^ ~\a[22] ) | (~\a[20]  ^ ~\a[21] )) & (new_n164_ | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ))));
  assign new_n403_ = ((new_n393_ | (new_n387_ & ~new_n388_) | (~new_n387_ & new_n388_)) & ((~new_n394_ & ~new_n396_) | (~new_n393_ & (~new_n387_ | new_n388_) & (new_n387_ | ~new_n388_)) | (new_n393_ & (~new_n387_ ^ ~new_n388_)))) ^ (new_n402_ ^ (new_n390_ ^ (new_n384_ | (new_n387_ & ~new_n388_))));
  assign new_n404_ = new_n397_ ^ (new_n394_ | new_n396_);
  assign new_n405_ = (~new_n403_ ^ \a[20] ) ^ ((~new_n404_ | ~\a[20] ) & ((new_n404_ & \a[20] ) | (~new_n404_ & ~\a[20] ) | ((~new_n166_ | ~\a[20] ) & (new_n154_ | (new_n166_ & \a[20] ) | (~new_n166_ & ~\a[20] )))));
  assign new_n406_ = ((new_n166_ & \a[20] ) | (~new_n154_ & (new_n166_ | \a[20] ) & (~new_n166_ | ~\a[20] ))) ^ (~new_n404_ ^ ~\a[20] );
  assign new_n407_ = (~\a[17]  | (new_n154_ & ~new_n165_) | (~new_n154_ & new_n165_)) & (((~new_n174_ | ~\a[17] ) & ((new_n174_ & \a[17] ) | (~new_n174_ & ~\a[17] ) | ((~new_n54_ | ~\a[17] ) & ((new_n54_ & \a[17] ) | (~new_n54_ & ~\a[17] ) | (~new_n176_ & (new_n177_ | ~new_n220_)))))) | (\a[17]  & (~new_n154_ | new_n165_) & (new_n154_ | ~new_n165_)) | (~\a[17]  & (~new_n154_ ^ ~new_n165_)));
  assign new_n408_ = \a[17]  ^ ((new_n404_ ^ \a[20] ) ^ ((new_n166_ & \a[20] ) | (~new_n154_ & (new_n166_ | \a[20] ) & (~new_n166_ | ~\a[20] ))));
  assign new_n409_ = (new_n405_ ^ \a[17] ) ^ ((~new_n407_ & new_n408_) | (new_n406_ & \a[17] ));
  assign new_n410_ = \a[14]  & (~new_n407_ | new_n408_) & (new_n407_ | ~new_n408_);
  assign new_n411_ = (~new_n153_ | ~\a[14] ) & ((new_n153_ & \a[14] ) | (~new_n153_ & ~\a[14] ) | ((~new_n221_ | ~\a[14] ) & ((new_n221_ & \a[14] ) | (~new_n221_ & ~\a[14] ) | ((~\a[14]  | (new_n53_ & (new_n176_ | (~new_n177_ & new_n220_))) | (~new_n53_ & ~new_n176_ & (new_n177_ | ~new_n220_))) & (((~\a[14]  | (~new_n177_ & new_n220_) | (new_n177_ & ~new_n220_)) & (new_n222_ | (\a[14]  & (new_n177_ | ~new_n220_) & (~new_n177_ | new_n220_)) | (~\a[14]  & (new_n177_ ^ new_n220_)))) | (\a[14]  & (~new_n53_ | (~new_n176_ & (new_n177_ | ~new_n220_))) & (new_n53_ | new_n176_ | (~new_n177_ & new_n220_))) | (~\a[14]  & (~new_n53_ ^ (new_n176_ | (~new_n177_ & new_n220_)))))))));
  assign new_n412_ = \a[14]  ^ (new_n407_ ^ ~new_n408_);
  assign new_n413_ = (~new_n414_ ^ ~\a[17] ) ^ ((new_n381_ & \a[17] ) | ((~new_n381_ | ~\a[17] ) & (new_n381_ | \a[17] ) & ((new_n405_ & \a[17] ) | ((~new_n405_ | ~\a[17] ) & (new_n405_ | \a[17] ) & ((~new_n407_ & new_n408_) | (new_n406_ & \a[17] ))))));
  assign new_n414_ = (~\a[20]  ^ (new_n415_ ^ ~new_n417_)) ^ ((~new_n382_ | ~\a[20] ) & ((new_n382_ & \a[20] ) | (~new_n382_ & ~\a[20] ) | ((~new_n403_ | ~\a[20] ) & ((new_n403_ & \a[20] ) | (~new_n403_ & ~\a[20] ) | ((~new_n404_ | ~\a[20] ) & ((new_n404_ & \a[20] ) | (~new_n404_ & ~\a[20] ) | ((~new_n166_ | ~\a[20] ) & (new_n154_ | (new_n166_ & \a[20] ) | (~new_n166_ & ~\a[20] )))))))));
  assign new_n415_ = (~new_n416_ | ~\a[23] ) & ((new_n416_ & \a[23] ) | (~new_n416_ & ~\a[23] ) | ((~new_n383_ | new_n402_) & ((new_n383_ & ~new_n402_) | (~new_n383_ & new_n402_) | (~new_n392_ & (~new_n397_ | (~new_n394_ & ~new_n396_))))));
  assign new_n416_ = new_n400_ ^ (new_n399_ | (new_n390_ & (new_n384_ | (new_n387_ & ~new_n388_))));
  assign new_n417_ = \a[23]  ^ (new_n420_ ^ (new_n419_ | (~new_n418_ & new_n400_)));
  assign new_n418_ = ~new_n399_ & (~new_n390_ | (~new_n384_ & (~new_n387_ | new_n388_)));
  assign new_n419_ = (new_n401_ ^ ~\a[26] ) & ((\b[11]  & (\a[26]  ^ \a[27] )) | (\b[10]  & \a[27]  & (\a[26]  | ~\a[27] ) & (~\a[26]  | \a[27] )));
  assign new_n420_ = ~new_n422_ ^ (new_n421_ ^ ~\a[26] );
  assign new_n421_ = ((\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (~\b[14]  ^ ((\b[13]  & \b[14] ) | (~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] ))))) & (~\b[13]  | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (~\a[24]  ^ ~\a[25] ) | (~\a[23]  ^ ~\a[24] )) & (~\b[14]  | (~\a[24]  & ~\a[25] ) | (\a[24]  & \a[25] ) | (~\a[23]  ^ ~\a[24] ));
  assign new_n422_ = (~\b[11]  | ~\a[27]  | (\a[26]  & ~\a[27] ) | (~\a[26]  & \a[27] )) & (~\b[12]  | (\a[26]  ^ ~\a[27] ));
  assign new_n423_ = (new_n380_ ^ \a[14] ) ^ ((new_n409_ & \a[14] ) | ((~new_n409_ | ~\a[14] ) & (new_n409_ | \a[14] ) & (new_n410_ | (~new_n411_ & new_n412_))));
  assign new_n424_ = (new_n410_ | (~new_n411_ & new_n412_)) ^ (new_n409_ ^ \a[14] );
  assign new_n425_ = new_n411_ ^ ~new_n412_;
  assign new_n426_ = (~new_n52_ | ~\a[11] ) & ((new_n52_ & \a[11] ) | (~new_n52_ & ~\a[11] ) | ((~new_n269_ | ~\a[11] ) & ((new_n269_ & \a[11] ) | (~new_n269_ & ~\a[11] ) | ((~\a[11]  | (new_n270_ & ~new_n320_) | (~new_n270_ & new_n320_)) & (new_n271_ | (\a[11]  & (~new_n270_ | new_n320_) & (new_n270_ | ~new_n320_)) | (~\a[11]  & (~new_n270_ ^ ~new_n320_)))))));
  assign new_n427_ = \a[8]  ^ (new_n428_ ^ ~new_n440_);
  assign new_n428_ = (~\a[11]  | (~new_n429_ & new_n430_) | (new_n429_ & ~new_n430_)) & ((\a[11]  & (new_n429_ | ~new_n430_) & (~new_n429_ | new_n430_)) | (~\a[11]  & (new_n429_ ^ new_n430_)) | ((~new_n379_ | ~\a[11] ) & ((new_n379_ & \a[11] ) | (~new_n379_ & ~\a[11] ) | ((~new_n423_ | ~\a[11] ) & ((new_n423_ & \a[11] ) | (~new_n423_ & ~\a[11] ) | ((~new_n424_ | ~\a[11] ) & ((new_n424_ & \a[11] ) | (~new_n424_ & ~\a[11] ) | ((~new_n425_ | ~\a[11] ) & (new_n426_ | (new_n425_ & \a[11] ) | (~new_n425_ & ~\a[11] ))))))))));
  assign new_n429_ = (~new_n413_ | ~\a[14] ) & ((new_n413_ & \a[14] ) | (~new_n413_ & ~\a[14] ) | ((~new_n380_ | ~\a[14] ) & ((~new_n380_ & ~\a[14] ) | (new_n380_ & \a[14] ) | ((~new_n409_ | ~\a[14] ) & ((~new_n410_ & (new_n411_ | ~new_n412_)) | (new_n409_ & \a[14] ) | (~new_n409_ & ~\a[14] ))))));
  assign new_n430_ = ~new_n431_ ^ ~\a[14] ;
  assign new_n431_ = (\a[17]  ^ (new_n432_ ^ ~new_n433_)) ^ ((new_n414_ & \a[17] ) | ((~new_n414_ | ~\a[17] ) & (new_n414_ | \a[17] ) & ((new_n381_ & \a[17] ) | ((~new_n381_ | ~\a[17] ) & (new_n381_ | \a[17] ) & ((new_n405_ & \a[17] ) | ((~new_n405_ | ~\a[17] ) & (new_n405_ | \a[17] ) & ((new_n406_ & \a[17] ) | (~new_n407_ & (~new_n406_ | ~\a[17] ) & (new_n406_ | \a[17] )))))))));
  assign new_n432_ = (~\a[20]  | (new_n415_ & ~new_n417_) | (~new_n415_ & new_n417_)) & ((\a[20]  & (~new_n415_ | new_n417_) & (new_n415_ | ~new_n417_)) | (~\a[20]  & (~new_n415_ ^ ~new_n417_)) | ((~new_n382_ | ~\a[20] ) & ((new_n382_ & \a[20] ) | (~new_n382_ & ~\a[20] ) | ((~new_n403_ | ~\a[20] ) & ((new_n403_ & \a[20] ) | (~new_n403_ & ~\a[20] ) | ((~new_n404_ | ~\a[20] ) & ((new_n404_ & \a[20] ) | (~new_n404_ & ~\a[20] ) | ((~new_n166_ | ~\a[20] ) & (new_n154_ | (new_n166_ & \a[20] ) | (~new_n166_ & ~\a[20] ))))))))));
  assign new_n433_ = \a[20]  ^ ((~\a[23]  ^ (~new_n435_ ^ new_n438_)) ^ ((~new_n434_ | ~\a[23] ) & (new_n415_ | (new_n434_ & \a[23] ) | (~new_n434_ & ~\a[23] ))));
  assign new_n434_ = new_n420_ ^ (new_n419_ | (~new_n418_ & new_n400_));
  assign new_n435_ = ~new_n436_ & ~new_n437_;
  assign new_n436_ = new_n420_ & (new_n419_ | (new_n400_ & (new_n399_ | (new_n390_ & (new_n384_ | (new_n387_ & ~new_n388_))))));
  assign new_n437_ = ~new_n422_ & (new_n421_ ^ ~\a[26] );
  assign new_n438_ = ((\b[13]  & (~\a[26]  ^ ~\a[27] )) | (\b[12]  & \a[27]  & (~\a[26]  | \a[27] ) & (\a[26]  | ~\a[27] ))) ^ (~\a[26]  ^ (~\b[14]  | (~new_n439_ & (~new_n59_ | ((~\b[13]  | ~\b[14] ) & (new_n114_ | (\b[13]  & \b[14] ) | (~\b[13]  & ~\b[14] )))))));
  assign new_n439_ = (\a[25]  | \a[26] ) & (~\a[25]  | ~\a[26] ) & (\a[23]  ^ ~\a[24] ) & (\a[24]  ^ ~\a[25] );
  assign new_n440_ = \a[11]  ^ (new_n441_ ^ ~new_n442_);
  assign new_n441_ = (~new_n431_ | ~\a[14] ) & ((new_n431_ & \a[14] ) | (~new_n431_ & ~\a[14] ) | ((~new_n413_ | ~\a[14] ) & ((new_n413_ & \a[14] ) | (~new_n413_ & ~\a[14] ) | ((~new_n380_ | ~\a[14] ) & ((new_n380_ & \a[14] ) | (~new_n380_ & ~\a[14] ) | ((~new_n409_ | ~\a[14] ) & ((new_n409_ & \a[14] ) | (~new_n409_ & ~\a[14] ) | (~new_n410_ & (new_n411_ | ~new_n412_)))))))));
  assign new_n442_ = ~\a[14]  ^ (~new_n445_ ^ ((new_n443_ & \a[17] ) | (~new_n444_ & (~new_n443_ | ~\a[17] ) & (new_n443_ | \a[17] ))));
  assign new_n443_ = new_n432_ ^ ~new_n433_;
  assign new_n444_ = (~new_n414_ | ~\a[17] ) & ((~new_n414_ & ~\a[17] ) | (new_n414_ & \a[17] ) | ((~new_n381_ | ~\a[17] ) & ((new_n381_ & \a[17] ) | (~new_n381_ & ~\a[17] ) | ((~new_n405_ | ~\a[17] ) & ((new_n405_ & \a[17] ) | (~new_n405_ & ~\a[17] ) | ((new_n407_ | ~new_n408_) & (~new_n406_ | ~\a[17] )))))));
  assign new_n445_ = ~\a[17]  ^ ((new_n447_ ^ ~\a[20] ) ^ ((new_n446_ & \a[20] ) | (~new_n432_ & (~new_n446_ | ~\a[20] ) & (new_n446_ | \a[20] ))));
  assign new_n446_ = ((~new_n434_ | ~\a[23] ) & (new_n415_ | (new_n434_ & \a[23] ) | (~new_n434_ & ~\a[23] ))) ^ (~\a[23]  ^ (~new_n435_ ^ new_n438_));
  assign new_n447_ = ~new_n448_ ^ ((~\a[23]  | (new_n435_ & ~new_n438_) | (~new_n435_ & new_n438_)) & (((~new_n434_ | ~\a[23] ) & (new_n415_ | (new_n434_ & \a[23] ) | (~new_n434_ & ~\a[23] ))) | (\a[23]  & (~new_n435_ | new_n438_) & (new_n435_ | ~new_n438_)) | (~\a[23]  & (~new_n435_ ^ ~new_n438_))));
  assign new_n448_ = \a[23]  ^ (new_n450_ ^ (new_n449_ | (new_n438_ & (new_n436_ | new_n437_))));
  assign new_n449_ = ((\b[13]  & (~\a[26]  ^ ~\a[27] )) | (\b[12]  & \a[27]  & (~\a[26]  | \a[27] ) & (\a[26]  | ~\a[27] ))) & (~\a[26]  ^ (~\b[14]  | (~new_n439_ & (~new_n59_ | ((~\b[13]  | ~\b[14] ) & (new_n114_ | (\b[13]  & \b[14] ) | (~\b[13]  & ~\b[14] )))))));
  assign new_n450_ = \a[26]  ? ((~\a[27]  | ~\b[13] ) & (~\b[14]  | (\a[26]  ^ ~\a[27] ))) : (\a[27]  & \b[14] );
  assign new_n451_ = ((\a[8]  & ((new_n423_ & \a[11] ) | (~new_n423_ & ~\a[11] ) | ((~new_n424_ | ~\a[11] ) & ((new_n424_ & \a[11] ) | (~new_n424_ & ~\a[11] ) | ((~new_n425_ | ~\a[11] ) & (new_n426_ | (new_n425_ & \a[11] ) | (~new_n425_ & ~\a[11] )))))) & ((new_n423_ ^ \a[11] ) | (new_n424_ & \a[11] ) | ((~new_n424_ | ~\a[11] ) & (new_n424_ | \a[11] ) & ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] )))))) | ((~\a[8]  | ((~new_n423_ | ~\a[11] ) & (new_n423_ | \a[11] ) & ((new_n424_ & \a[11] ) | ((~new_n424_ | ~\a[11] ) & (new_n424_ | \a[11] ) & ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] )))))) | ((~new_n423_ ^ \a[11] ) & (~new_n424_ | ~\a[11] ) & ((new_n424_ & \a[11] ) | (~new_n424_ & ~\a[11] ) | ((~new_n425_ | ~\a[11] ) & (new_n426_ | (new_n425_ & \a[11] ) | (~new_n425_ & ~\a[11] )))))) & (\a[8]  | ((new_n423_ ^ \a[11] ) ^ ((new_n424_ & \a[11] ) | ((~new_n424_ | ~\a[11] ) & (new_n424_ | \a[11] ) & ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] ))))))) & ((\a[8]  & ((new_n424_ & \a[11] ) | (~new_n424_ & ~\a[11] ) | ((~new_n425_ | ~\a[11] ) & (new_n426_ | (new_n425_ & \a[11] ) | (~new_n425_ & ~\a[11] )))) & ((new_n424_ ^ \a[11] ) | (new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] )))) | ((~\a[8]  | ((~new_n424_ | ~\a[11] ) & (new_n424_ | \a[11] ) & ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] )))) | ((~new_n424_ ^ \a[11] ) & (~new_n425_ | ~\a[11] ) & (new_n426_ | (new_n425_ & \a[11] ) | (~new_n425_ & ~\a[11] )))) & (\a[8]  | ((new_n424_ ^ \a[11] ) ^ ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] ))))) & ((\a[8]  & (new_n426_ | (new_n425_ & \a[11] ) | (~new_n425_ & ~\a[11] )) & (~new_n426_ | (new_n425_ ^ \a[11] ))) | (~new_n50_ & (~\a[8]  | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] )) | (new_n426_ & (~new_n425_ ^ \a[11] ))) & (\a[8]  | (~new_n426_ ^ (new_n425_ ^ \a[11] ))))))))) ^ (\a[8]  ^ ((new_n379_ ^ \a[11] ) ^ ((new_n423_ & \a[11] ) | ((~new_n423_ | ~\a[11] ) & (new_n423_ | \a[11] ) & ((new_n424_ & \a[11] ) | ((~new_n424_ | ~\a[11] ) & (new_n424_ | \a[11] ) & ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] )))))))));
  assign new_n452_ = (~\a[5]  | (new_n453_ & ~new_n457_) | (~new_n453_ & new_n457_)) & ((\a[5]  & (~new_n453_ | new_n457_) & (new_n453_ | ~new_n457_)) | (~\a[5]  & (~new_n453_ ^ ~new_n457_)) | ((~new_n458_ | ~\a[5] ) & ((new_n458_ & \a[5] ) | (~new_n458_ & ~\a[5] ) | ((~new_n459_ | ~\a[5] ) & ((new_n459_ & \a[5] ) | (~new_n459_ & ~\a[5] ) | ((~new_n460_ | ~\a[5] ) & ((new_n460_ & \a[5] ) | (~new_n460_ & ~\a[5] ) | ((~new_n461_ | ~\a[5] ) & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] ))))))))));
  assign new_n453_ = (~\a[8]  | (new_n454_ & ~new_n455_) | (~new_n454_ & new_n455_)) & (((~new_n456_ | ~\a[8] ) & ((new_n456_ & \a[8] ) | (~new_n456_ & ~\a[8] ) | ((~new_n51_ | ~\a[8] ) & ((new_n51_ & \a[8] ) | (~new_n51_ & ~\a[8] ) | (~new_n321_ & (new_n322_ | ~new_n378_)))))) | (\a[8]  & (~new_n454_ | new_n455_) & (new_n454_ | ~new_n455_)) | (~\a[8]  & (~new_n454_ ^ ~new_n455_)));
  assign new_n454_ = (~\a[11]  | (new_n411_ & ~new_n412_) | (~new_n411_ & new_n412_)) & ((\a[11]  & (~new_n411_ | new_n412_) & (new_n411_ | ~new_n412_)) | (~\a[11]  & (~new_n411_ ^ ~new_n412_)) | ((~new_n52_ | ~\a[11] ) & ((new_n52_ & \a[11] ) | (~new_n52_ & ~\a[11] ) | ((~new_n269_ | ~\a[11] ) & ((new_n269_ & \a[11] ) | (~new_n269_ & ~\a[11] ) | ((~\a[11]  | (~new_n270_ & new_n320_) | (new_n270_ & ~new_n320_)) & (new_n271_ | (\a[11]  & (new_n270_ | ~new_n320_) & (~new_n270_ | new_n320_)) | (~\a[11]  & (new_n270_ ^ new_n320_)))))))));
  assign new_n455_ = \a[11]  ^ ((new_n410_ | (~new_n411_ & new_n412_)) ^ (new_n409_ ^ \a[14] ));
  assign new_n456_ = (\a[11]  ^ (new_n411_ ^ ~new_n412_)) ^ ((new_n52_ & \a[11] ) | ((~new_n52_ | ~\a[11] ) & (new_n52_ | \a[11] ) & ((new_n269_ & \a[11] ) | ((~new_n269_ | ~\a[11] ) & (new_n269_ | \a[11] ) & ((\a[11]  & (new_n270_ | ~new_n320_) & (~new_n270_ | new_n320_)) | (~new_n271_ & (~\a[11]  | (~new_n270_ & new_n320_) | (new_n270_ & ~new_n320_)) & (\a[11]  | (~new_n270_ ^ new_n320_))))))));
  assign new_n457_ = \a[8]  ^ ((new_n423_ ^ \a[11] ) ^ ((new_n424_ & \a[11] ) | ((~new_n424_ | ~\a[11] ) & (new_n424_ | \a[11] ) & ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] ))))));
  assign new_n458_ = ((new_n456_ & \a[8] ) | ((~new_n456_ | ~\a[8] ) & (new_n456_ | \a[8] ) & ((new_n51_ & \a[8] ) | ((~new_n51_ | ~\a[8] ) & (new_n51_ | \a[8] ) & (new_n321_ | (~new_n322_ & new_n378_)))))) ^ (\a[8]  ^ (new_n454_ ^ ~new_n455_));
  assign new_n459_ = (new_n456_ ^ \a[8] ) ^ ((new_n51_ & \a[8] ) | ((~new_n51_ | ~\a[8] ) & (new_n51_ | \a[8] ) & (new_n321_ | (~new_n322_ & new_n378_))));
  assign new_n460_ = (new_n321_ | (~new_n322_ & new_n378_)) ^ (new_n51_ ^ \a[8] );
  assign new_n461_ = new_n322_ ^ ~new_n378_;
  assign new_n462_ = (~new_n463_ | ~\a[5] ) & ((~new_n463_ & ~\a[5] ) | (new_n463_ & \a[5] ) | ((~\a[5]  | ((~new_n324_ | ~\a[8] ) & (new_n324_ | \a[8] ) & ((new_n325_ & \a[8] ) | ((~new_n325_ | ~\a[8] ) & (new_n325_ | \a[8] ) & ((new_n326_ & \a[8] ) | (~new_n328_ & (~new_n326_ | ~\a[8] ) & (new_n326_ | \a[8] )))))) | ((~new_n324_ ^ \a[8] ) & (~new_n325_ | ~\a[8] ) & ((new_n325_ & \a[8] ) | (~new_n325_ & ~\a[8] ) | ((~new_n326_ | ~\a[8] ) & (new_n328_ | (new_n326_ & \a[8] ) | (~new_n326_ & ~\a[8] )))))) & ((\a[5]  & ((new_n324_ & \a[8] ) | (~new_n324_ & ~\a[8] ) | ((~new_n325_ | ~\a[8] ) & ((new_n325_ & \a[8] ) | (~new_n325_ & ~\a[8] ) | ((~new_n326_ | ~\a[8] ) & (new_n328_ | (new_n326_ & \a[8] ) | (~new_n326_ & ~\a[8] )))))) & ((new_n324_ ^ \a[8] ) | (new_n325_ & \a[8] ) | ((~new_n325_ | ~\a[8] ) & (new_n325_ | \a[8] ) & ((new_n326_ & \a[8] ) | (~new_n328_ & (~new_n326_ | ~\a[8] ) & (new_n326_ | \a[8] )))))) | (~\a[5]  & ((~new_n324_ ^ \a[8] ) ^ ((new_n325_ & \a[8] ) | ((~new_n325_ | ~\a[8] ) & (new_n325_ | \a[8] ) & ((new_n326_ & \a[8] ) | (~new_n328_ & (~new_n326_ | ~\a[8] ) & (new_n326_ | \a[8] ))))))) | ((~\a[5]  | ((~new_n325_ | ~\a[8] ) & (new_n325_ | \a[8] ) & ((new_n326_ & \a[8] ) | (~new_n328_ & (~new_n326_ | ~\a[8] ) & (new_n326_ | \a[8] )))) | ((~new_n325_ ^ \a[8] ) & (~new_n326_ | ~\a[8] ) & (new_n328_ | (new_n326_ & \a[8] ) | (~new_n326_ & ~\a[8] )))) & (new_n464_ | (\a[5]  & ((new_n325_ & \a[8] ) | (~new_n325_ & ~\a[8] ) | ((~new_n326_ | ~\a[8] ) & (new_n328_ | (new_n326_ & \a[8] ) | (~new_n326_ & ~\a[8] )))) & ((new_n325_ ^ \a[8] ) | (new_n326_ & \a[8] ) | (~new_n328_ & (~new_n326_ | ~\a[8] ) & (new_n326_ | \a[8] )))) | (~\a[5]  & ((~new_n325_ ^ \a[8] ) ^ ((new_n326_ & \a[8] ) | (~new_n328_ & (~new_n326_ | ~\a[8] ) & (new_n326_ | \a[8] ))))))))));
  assign new_n463_ = ((new_n324_ & \a[8] ) | ((~new_n324_ | ~\a[8] ) & (new_n324_ | \a[8] ) & ((new_n325_ & \a[8] ) | (((new_n326_ & \a[8] ) | (~new_n328_ & (new_n326_ | \a[8] ) & (~new_n326_ | ~\a[8] ))) & (~new_n325_ | ~\a[8] ) & (new_n325_ | \a[8] ))))) ^ (\a[8]  ^ (new_n271_ ^ ~new_n323_));
  assign new_n464_ = (~\a[5]  | (new_n328_ & ~new_n465_) | (~new_n328_ & new_n465_)) & (((~new_n466_ | ~\a[5] ) & ((new_n466_ & \a[5] ) | (~new_n466_ & ~\a[5] ) | ((~new_n467_ | ~\a[5] ) & (((~new_n468_ | ~\a[5] ) & (new_n470_ | (~new_n468_ & ~\a[5] ) | (new_n468_ & \a[5] ))) | (new_n467_ & \a[5] ) | (~new_n467_ & ~\a[5] ))))) | (\a[5]  & (~new_n328_ | new_n465_) & (new_n328_ | ~new_n465_)) | (~\a[5]  & (~new_n328_ ^ ~new_n465_)));
  assign new_n465_ = \a[8]  ^ (new_n273_ ^ ~new_n327_);
  assign new_n466_ = (new_n330_ ^ \a[8] ) ^ ((\a[8]  & (((~new_n276_ | ~\a[11] ) & ((new_n276_ & \a[11] ) | (~new_n276_ & ~\a[11] ) | ((~new_n277_ | ~\a[11] ) & (new_n279_ | (new_n277_ & \a[11] ) | (~new_n277_ & ~\a[11] ))))) | (new_n329_ & \a[11] ) | (~new_n329_ & ~\a[11] )) & ((new_n276_ & \a[11] ) | ((~new_n276_ | ~\a[11] ) & (new_n276_ | \a[11] ) & ((new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] )))) | (new_n329_ ^ \a[11] ))) | ((~\a[8]  | (((new_n276_ & \a[11] ) | ((~new_n276_ | ~\a[11] ) & (new_n276_ | \a[11] ) & ((new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] ))))) & (~new_n329_ | ~\a[11] ) & (new_n329_ | \a[11] )) | ((~new_n276_ | ~\a[11] ) & ((new_n276_ & \a[11] ) | (~new_n276_ & ~\a[11] ) | ((~new_n277_ | ~\a[11] ) & (new_n279_ | (new_n277_ & \a[11] ) | (~new_n277_ & ~\a[11] )))) & (~new_n329_ ^ \a[11] ))) & (\a[8]  | (((new_n276_ & \a[11] ) | ((~new_n276_ | ~\a[11] ) & (new_n276_ | \a[11] ) & ((new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] ))))) ^ (new_n329_ ^ \a[11] ))) & ((\a[8]  & ((new_n276_ & \a[11] ) | (~new_n276_ & ~\a[11] ) | ((~new_n277_ | ~\a[11] ) & (new_n279_ | (new_n277_ & \a[11] ) | (~new_n277_ & ~\a[11] )))) & ((new_n276_ ^ \a[11] ) | (new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] )))) | (~new_n331_ & (~\a[8]  | ((~new_n276_ | ~\a[11] ) & (new_n276_ | \a[11] ) & ((new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] )))) | ((~new_n276_ ^ \a[11] ) & (~new_n277_ | ~\a[11] ) & (new_n279_ | (new_n277_ & \a[11] ) | (~new_n277_ & ~\a[11] )))) & (\a[8]  | ((new_n276_ ^ \a[11] ) ^ ((new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] )))))))));
  assign new_n467_ = (\a[8]  ^ ((~new_n329_ ^ ~\a[11] ) ^ ((new_n276_ & \a[11] ) | ((~new_n276_ | ~\a[11] ) & (new_n276_ | \a[11] ) & ((new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] ))))))) ^ ((\a[8]  & ((new_n276_ & \a[11] ) | (~new_n276_ & ~\a[11] ) | ((~new_n277_ | ~\a[11] ) & (new_n279_ | (new_n277_ & \a[11] ) | (~new_n277_ & ~\a[11] )))) & ((new_n276_ ^ \a[11] ) | (new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] )))) | (~new_n331_ & (~\a[8]  | ((~new_n276_ | ~\a[11] ) & (new_n276_ | \a[11] ) & ((new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] )))) | ((~new_n276_ ^ \a[11] ) & (~new_n277_ | ~\a[11] ) & (new_n279_ | (new_n277_ & \a[11] ) | (~new_n277_ & ~\a[11] )))) & (\a[8]  | ((new_n276_ ^ \a[11] ) ^ ((new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] )))))));
  assign new_n468_ = new_n469_ ^ ~new_n331_;
  assign new_n469_ = \a[8]  ^ ((new_n276_ ^ \a[11] ) ^ ((new_n277_ & \a[11] ) | (~new_n279_ & (~new_n277_ | ~\a[11] ) & (new_n277_ | \a[11] ))));
  assign new_n470_ = (~new_n472_ | ~\a[5] ) & ((new_n472_ & \a[5] ) | (~new_n472_ & ~\a[5] ) | ((~\a[5]  | (((new_n334_ & \a[8] ) | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] ))))) & (~new_n471_ | ~\a[8] ) & (new_n471_ | \a[8] )) | ((~new_n334_ | ~\a[8] ) & ((new_n334_ & \a[8] ) | (~new_n334_ & ~\a[8] ) | ((~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))) & (~new_n471_ ^ \a[8] ))) & ((\a[5]  & (((~new_n334_ | ~\a[8] ) & ((new_n334_ & \a[8] ) | (~new_n334_ & ~\a[8] ) | ((~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] ))))) | (new_n471_ & \a[8] ) | (~new_n471_ & ~\a[8] )) & ((new_n334_ & \a[8] ) | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))) | (new_n471_ ^ \a[8] ))) | (~\a[5]  & (((~new_n334_ | ~\a[8] ) & ((new_n334_ & \a[8] ) | (~new_n334_ & ~\a[8] ) | ((~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] ))))) ^ (new_n471_ ^ \a[8] ))) | ((~\a[5]  | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))) | ((~new_n334_ ^ \a[8] ) & (~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))) & (new_n473_ | (\a[5]  & ((new_n334_ & \a[8] ) | (~new_n334_ & ~\a[8] ) | ((~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))) & ((new_n334_ ^ \a[8] ) | (new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))) | (~\a[5]  & ((~new_n334_ ^ \a[8] ) ^ ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] ))))))))));
  assign new_n471_ = ~new_n332_ ^ (~new_n280_ ^ new_n318_);
  assign new_n472_ = ((\a[8]  & (new_n332_ | (~new_n280_ & new_n318_) | (new_n280_ & ~new_n318_)) & (~new_n332_ | (~new_n280_ ^ new_n318_))) | (((new_n334_ & \a[8] ) | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] ))))) & (~\a[8]  | (~new_n332_ & (new_n280_ | ~new_n318_) & (~new_n280_ | new_n318_)) | (new_n332_ & (new_n280_ ^ new_n318_))) & (\a[8]  | (~new_n332_ ^ (~new_n280_ ^ new_n318_))))) ^ (\a[8]  ^ (new_n333_ ^ ((new_n280_ & ~new_n318_) | (~new_n332_ & (new_n280_ | ~new_n318_) & (~new_n280_ | new_n318_)))));
  assign new_n473_ = (~\a[5]  | (new_n337_ & ~new_n474_) | (~new_n337_ & new_n474_)) & (((~new_n475_ | ~\a[5] ) & ((new_n475_ & \a[5] ) | (~new_n475_ & ~\a[5] ) | ((~new_n477_ | ~\a[5] ) & (((~new_n478_ | ~\a[5] ) & (new_n480_ | (~new_n478_ & ~\a[5] ) | (new_n478_ & \a[5] ))) | (new_n477_ & \a[5] ) | (~new_n477_ & ~\a[5] ))))) | (\a[5]  & (~new_n337_ | new_n474_) & (new_n337_ | ~new_n474_)) | (~\a[5]  & (~new_n337_ ^ ~new_n474_)));
  assign new_n474_ = \a[8]  ^ (new_n283_ ^ ~new_n336_);
  assign new_n475_ = new_n476_ ^ (new_n339_ | (~new_n339_ & ~new_n375_ & ((~new_n377_ & (new_n291_ | ~new_n314_) & (~new_n291_ | new_n314_)) | (~new_n341_ & (new_n377_ | (~new_n291_ & new_n314_) | (new_n291_ & ~new_n314_)) & (~new_n377_ | (~new_n291_ ^ new_n314_))))));
  assign new_n476_ = ~new_n376_ ^ ((new_n286_ | (new_n315_ & (new_n288_ | (~new_n291_ & new_n314_)))) ^ (new_n284_ ^ ~new_n316_));
  assign new_n477_ = (~new_n339_ & ~new_n375_) ^ ((~new_n377_ & (~new_n291_ | new_n314_) & (new_n291_ | ~new_n314_)) | (~new_n341_ & (~new_n377_ | (new_n291_ ^ ~new_n314_)) & (new_n377_ | (new_n291_ & ~new_n314_) | (~new_n291_ & new_n314_))));
  assign new_n478_ = new_n341_ ^ ~new_n479_;
  assign new_n479_ = ~new_n377_ ^ (new_n291_ ^ ~new_n314_);
  assign new_n480_ = (~new_n481_ | new_n520_) & ((new_n481_ & ~new_n520_) | (~new_n481_ & new_n520_) | (~new_n482_ & (((new_n521_ | (~new_n349_ & new_n372_) | (new_n349_ & ~new_n372_)) & (new_n484_ | (~new_n521_ & (new_n349_ | ~new_n372_) & (~new_n349_ | new_n372_)) | (new_n521_ & (new_n349_ ^ new_n372_)))) | new_n482_ | new_n519_)));
  assign new_n481_ = (new_n344_ | (new_n373_ & (new_n346_ | (~new_n349_ & new_n372_)))) ^ (new_n342_ ^ ~new_n374_);
  assign new_n482_ = ~new_n483_ & (~new_n373_ | (~new_n346_ & (new_n349_ | ~new_n372_))) & (new_n373_ | new_n346_ | (~new_n349_ & new_n372_));
  assign new_n483_ = \a[5]  ^ (((\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\b[14]  ^ ((\b[13]  & \b[14] ) | (~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] ))))) & (~\b[14]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[13]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n484_ = (~new_n485_ | new_n518_) & ((~new_n487_ & (~new_n517_ | (~new_n489_ & (new_n492_ | ~new_n516_)))) | (new_n485_ & ~new_n518_) | (~new_n485_ & new_n518_));
  assign new_n485_ = new_n486_ ^ (new_n352_ | (new_n368_ & ((~new_n371_ & (new_n302_ | (~new_n301_ & new_n309_) | (new_n301_ & ~new_n309_)) & (~new_n302_ | (~new_n301_ ^ new_n309_))) | (~new_n354_ & (new_n371_ | (~new_n302_ & (new_n301_ | ~new_n309_) & (~new_n301_ | new_n309_)) | (new_n302_ & (new_n301_ ^ new_n309_))) & (~new_n371_ | (~new_n302_ ^ (~new_n301_ ^ new_n309_)))))));
  assign new_n486_ = ~new_n369_ ^ ((new_n297_ ^ ~new_n298_) ^ ((new_n299_ & ~new_n300_) | ((new_n299_ | ~new_n300_) & (~new_n299_ | new_n300_) & ((~new_n301_ & new_n309_) | (~new_n302_ & (new_n301_ | ~new_n309_) & (~new_n301_ | new_n309_))))));
  assign new_n487_ = ~new_n488_ & (~new_n368_ | ((new_n371_ | (~new_n302_ & (new_n301_ | ~new_n309_) & (~new_n301_ | new_n309_)) | (new_n302_ & (new_n301_ ^ new_n309_))) & (new_n354_ | (~new_n371_ & (new_n302_ | (~new_n301_ & new_n309_) | (new_n301_ & ~new_n309_)) & (~new_n302_ | (~new_n301_ ^ new_n309_))) | (new_n371_ & (new_n302_ ^ (~new_n301_ ^ new_n309_)))))) & (new_n368_ | (~new_n371_ & (new_n302_ | (~new_n301_ & new_n309_) | (new_n301_ & ~new_n309_)) & (~new_n302_ | (~new_n301_ ^ new_n309_))) | (~new_n354_ & (new_n371_ | (~new_n302_ & (new_n301_ | ~new_n309_) & (~new_n301_ | new_n309_)) | (new_n302_ & (new_n301_ ^ new_n309_))) & (~new_n371_ | (~new_n302_ ^ (~new_n301_ ^ new_n309_)))));
  assign new_n488_ = \a[5]  ^ ((~new_n106_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[11]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[12]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[10]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n489_ = ~new_n491_ & (~new_n354_ | new_n490_) & (new_n354_ | ~new_n490_);
  assign new_n490_ = ~new_n371_ ^ (~new_n302_ ^ (new_n301_ ^ ~new_n309_));
  assign new_n491_ = \a[5]  ^ ((~new_n112_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[10]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[11]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[9]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n492_ = (~new_n494_ | new_n513_) & ((new_n494_ & ~new_n513_) | (~new_n494_ & new_n513_) | (~new_n495_ & (~new_n497_ | ((new_n515_ | (new_n493_ & ~new_n360_) | (~new_n493_ & new_n360_)) & (new_n498_ | (~new_n515_ & (~new_n493_ | new_n360_) & (new_n493_ | ~new_n360_)) | (new_n515_ & (~new_n493_ ^ ~new_n360_)))))));
  assign new_n493_ = new_n359_ ^ ~new_n367_;
  assign new_n494_ = (new_n355_ ^ ~new_n356_) ^ ((new_n357_ & ~new_n358_) | ((new_n357_ | ~new_n358_) & (~new_n357_ | new_n358_) & ((~new_n359_ & new_n367_) | (~new_n360_ & (new_n359_ | ~new_n367_) & (~new_n359_ | new_n367_)))));
  assign new_n495_ = ~new_n496_ & ((new_n357_ & ~new_n358_) | (~new_n357_ & new_n358_) | ((new_n359_ | ~new_n367_) & (new_n360_ | (~new_n359_ & new_n367_) | (new_n359_ & ~new_n367_)))) & ((new_n357_ ^ ~new_n358_) | (~new_n359_ & new_n367_) | (~new_n360_ & (new_n359_ | ~new_n367_) & (~new_n359_ | new_n367_)));
  assign new_n496_ = \a[5]  ^ (((\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[9]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[7]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n497_ = ~new_n496_ ^ ((new_n357_ ^ ~new_n358_) ^ ((~new_n359_ & new_n367_) | (~new_n360_ & (new_n359_ | ~new_n367_) & (~new_n359_ | new_n367_))));
  assign new_n498_ = (~new_n499_ | new_n500_) & ((new_n499_ & ~new_n500_) | (~new_n499_ & new_n500_) | ((~new_n501_ | new_n502_) & ((~new_n501_ & new_n502_) | (new_n501_ & ~new_n502_) | ((new_n503_ | ~new_n512_) & (new_n506_ | (~new_n503_ & new_n512_) | (new_n503_ & ~new_n512_))))));
  assign new_n499_ = (new_n364_ | (~new_n365_ & new_n366_)) ^ (new_n363_ ^ (~\a[8]  ^ (new_n362_ & (~new_n66_ | ~new_n361_))));
  assign new_n500_ = \a[5]  ^ ((~new_n75_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[6]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[7]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[5]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n501_ = new_n365_ ^ ~new_n366_;
  assign new_n502_ = \a[5]  ^ ((~new_n60_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[5]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[6]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[4]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n503_ = \a[5]  ^ (new_n505_ & (~new_n63_ | ~new_n504_));
  assign new_n504_ = (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (\a[4]  | \a[5] ) & (~\a[4]  | ~\a[5] );
  assign new_n505_ = (~\b[4]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[5]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[3]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n506_ = (~new_n508_ | (\a[5]  ^ (new_n507_ & (~new_n66_ | ~new_n504_)))) & ((~new_n509_ & (new_n510_ | ~new_n511_)) | (new_n508_ & (~\a[5]  ^ (new_n507_ & (~new_n66_ | ~new_n504_)))) | (~new_n508_ & (~\a[5]  | ~new_n507_ | (new_n66_ & new_n504_)) & (\a[5]  | (new_n507_ & (~new_n66_ | ~new_n504_)))));
  assign new_n507_ = (~\b[3]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[4]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[2]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n508_ = ((\b[0]  & (\a[5]  ^ ~\a[6] ) & (\a[6]  | \a[7] ) & (~\a[6]  | ~\a[7] )) | (\b[1]  & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (\a[7]  ^ ~\a[8] )) | ((\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[8]  & \b[0]  & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ));
  assign new_n509_ = \b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (~\b[0]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[1]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n510_ = \a[5]  ^ (((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[2]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )));
  assign new_n511_ = (\b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] )) ^ ((~\b[0]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[1]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )));
  assign new_n512_ = (~\a[8]  | ((~\b[0]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )))) ^ ((~\b[1]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[2]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )));
  assign new_n513_ = \a[5]  ^ (new_n514_ & (~new_n504_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n514_ = (~\b[9]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[10]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[8]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n515_ = \a[5]  ^ (((~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n80_ & (~\b[7]  ^ \b[8] )) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[7]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[8]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[6]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n516_ = ~new_n491_ ^ (new_n354_ ^ ~new_n490_);
  assign new_n517_ = ~new_n488_ ^ (new_n368_ ^ ((~new_n371_ & (new_n302_ | (~new_n301_ & new_n309_) | (new_n301_ & ~new_n309_)) & (~new_n302_ | (~new_n301_ ^ new_n309_))) | (~new_n354_ & (new_n371_ | (~new_n302_ & (new_n301_ | ~new_n309_) & (~new_n301_ | new_n309_)) | (new_n302_ & (new_n301_ ^ new_n309_))) & (~new_n371_ | (~new_n302_ ^ (~new_n301_ ^ new_n309_))))));
  assign new_n518_ = \a[5]  ^ ((~new_n149_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[12]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[13]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[11]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n519_ = new_n483_ & (~new_n373_ ^ (new_n346_ | (~new_n349_ & new_n372_)));
  assign new_n520_ = \a[5]  ^ (~\b[14]  | ((new_n164_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] ))));
  assign new_n521_ = \a[5]  ^ (((~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n114_ & (~\b[13]  ^ \b[14] )) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[13]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[14]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[12]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n522_ = (\a[11]  ^ (~new_n429_ ^ new_n430_)) ^ ((new_n379_ & \a[11] ) | ((~new_n379_ | ~\a[11] ) & (new_n379_ | \a[11] ) & ((new_n423_ & \a[11] ) | ((~new_n423_ | ~\a[11] ) & (new_n423_ | \a[11] ) & ((new_n424_ & \a[11] ) | ((~new_n424_ | ~\a[11] ) & (new_n424_ | \a[11] ) & ((new_n425_ & \a[11] ) | (~new_n426_ & (~new_n425_ | ~\a[11] ) & (new_n425_ | \a[11] )))))))));
  assign new_n523_ = \a[11]  ^ ((\a[14]  & (~new_n445_ | ((~new_n443_ | ~\a[17] ) & (new_n444_ | (new_n443_ & \a[17] ) | (~new_n443_ & ~\a[17] )))) & (new_n445_ | (new_n443_ & \a[17] ) | (~new_n444_ & (~new_n443_ | ~\a[17] ) & (new_n443_ | \a[17] )))) | (~new_n441_ & (~\a[14]  | (new_n445_ & ((new_n443_ & \a[17] ) | (~new_n444_ & (~new_n443_ | ~\a[17] ) & (new_n443_ | \a[17] )))) | (~new_n445_ & (~new_n443_ | ~\a[17] ) & (new_n444_ | (new_n443_ & \a[17] ) | (~new_n443_ & ~\a[17] )))) & (\a[14]  | (new_n445_ ^ ((new_n443_ & \a[17] ) | (~new_n444_ & (~new_n443_ | ~\a[17] ) & (new_n443_ | \a[17] )))))));
  assign new_n524_ = (~\a[20]  ^ ~\a[23] ) ^ (\a[8]  ^ ((\a[17]  & ((new_n447_ & \a[20] ) | (~new_n447_ & ~\a[20] ) | ((~new_n446_ | ~\a[20] ) & (new_n432_ | (new_n446_ & \a[20] ) | (~new_n446_ & ~\a[20] )))) & ((new_n447_ ^ \a[20] ) | (new_n446_ & \a[20] ) | (~new_n432_ & (~new_n446_ | ~\a[20] ) & (new_n446_ | \a[20] )))) | (((\a[17]  & (new_n432_ | (new_n446_ & \a[20] ) | (~new_n446_ & ~\a[20] )) & (~new_n432_ | (new_n446_ ^ \a[20] ))) | (~new_n444_ & (~\a[17]  | (~new_n432_ & (~new_n446_ | ~\a[20] ) & (new_n446_ | \a[20] )) | (new_n432_ & (~new_n446_ ^ \a[20] ))) & (\a[17]  | (~new_n432_ ^ (new_n446_ ^ \a[20] ))))) & (~\a[17]  | ((~new_n447_ | ~\a[20] ) & (new_n447_ | \a[20] ) & ((new_n446_ & \a[20] ) | (~new_n432_ & (~new_n446_ | ~\a[20] ) & (new_n446_ | \a[20] )))) | ((~new_n447_ ^ \a[20] ) & (~new_n446_ | ~\a[20] ) & (new_n432_ | (new_n446_ & \a[20] ) | (~new_n446_ & ~\a[20] )))) & (\a[17]  | ((new_n447_ ^ \a[20] ) ^ ((new_n446_ & \a[20] ) | (~new_n432_ & (~new_n446_ | ~\a[20] ) & (new_n446_ | \a[20] ))))))));
  assign new_n525_ = ((\a[5]  & (new_n49_ | (~new_n522_ & ~\a[8] ) | (new_n522_ & \a[8] )) & (~new_n49_ | (~new_n522_ ^ ~\a[8] ))) | (~new_n526_ & (~\a[5]  | (~new_n49_ & (new_n522_ | \a[8] ) & (~new_n522_ | ~\a[8] )) | (new_n49_ & (new_n522_ ^ ~\a[8] ))) & (\a[5]  | (~new_n49_ ^ (~new_n522_ ^ ~\a[8] ))))) ^ (\a[5]  ^ (new_n427_ ^ ((new_n522_ & \a[8] ) | (~new_n49_ & (new_n522_ | \a[8] ) & (~new_n522_ | ~\a[8] )))));
  assign new_n526_ = (~new_n451_ | ~\a[5] ) & (new_n452_ | (~new_n451_ & ~\a[5] ) | (new_n451_ & \a[5] ));
  assign new_n527_ = (~\a[2]  | (new_n526_ & ~new_n528_) | (~new_n526_ & new_n528_)) & (((~new_n529_ | ~\a[2] ) & (((~new_n588_ | ~\a[2] ) & (new_n530_ | (new_n588_ & \a[2] ) | (~new_n588_ & ~\a[2] ))) | (new_n529_ & \a[2] ) | (~new_n529_ & ~\a[2] ))) | (\a[2]  & (~new_n526_ | new_n528_) & (new_n526_ | ~new_n528_)) | (~\a[2]  & (~new_n526_ ^ ~new_n528_)));
  assign new_n528_ = \a[5]  ^ (~new_n49_ ^ (~new_n522_ ^ ~\a[8] ));
  assign new_n529_ = ~new_n452_ ^ (~new_n451_ ^ ~\a[5] );
  assign new_n530_ = (~\a[2]  | ((~new_n458_ | ~\a[5] ) & (new_n458_ | \a[5] ) & ((new_n459_ & \a[5] ) | ((~new_n459_ | ~\a[5] ) & (new_n459_ | \a[5] ) & ((new_n460_ & \a[5] ) | ((~new_n460_ | ~\a[5] ) & (new_n460_ | \a[5] ) & ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )))))))) | ((~new_n458_ ^ \a[5] ) & (~new_n459_ | ~\a[5] ) & ((new_n459_ & \a[5] ) | (~new_n459_ & ~\a[5] ) | ((~new_n460_ | ~\a[5] ) & ((new_n460_ & \a[5] ) | (~new_n460_ & ~\a[5] ) | ((~new_n461_ | ~\a[5] ) & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )))))))) & (((~\a[2]  | ((~new_n459_ | ~\a[5] ) & (new_n459_ | \a[5] ) & ((new_n460_ & \a[5] ) | ((~new_n460_ | ~\a[5] ) & (new_n460_ | \a[5] ) & ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )))))) | ((~new_n459_ ^ \a[5] ) & (~new_n460_ | ~\a[5] ) & ((new_n460_ & \a[5] ) | (~new_n460_ & ~\a[5] ) | ((~new_n461_ | ~\a[5] ) & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )))))) & ((\a[2]  & ((new_n459_ & \a[5] ) | (~new_n459_ & ~\a[5] ) | ((~new_n460_ | ~\a[5] ) & ((new_n460_ & \a[5] ) | (~new_n460_ & ~\a[5] ) | ((~new_n461_ | ~\a[5] ) & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )))))) & ((new_n459_ ^ \a[5] ) | (new_n460_ & \a[5] ) | ((~new_n460_ | ~\a[5] ) & (new_n460_ | \a[5] ) & ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )))))) | (~\a[2]  & ((~new_n459_ ^ \a[5] ) ^ ((new_n460_ & \a[5] ) | ((~new_n460_ | ~\a[5] ) & (new_n460_ | \a[5] ) & ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] ))))))) | ((~\a[2]  | ((~new_n460_ | ~\a[5] ) & (new_n460_ | \a[5] ) & ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )))) | ((~new_n460_ ^ \a[5] ) & (~new_n461_ | ~\a[5] ) & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )))) & ((\a[2]  & ((new_n460_ & \a[5] ) | (~new_n460_ & ~\a[5] ) | ((~new_n461_ | ~\a[5] ) & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )))) & ((new_n460_ ^ \a[5] ) | (new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )))) | (~\a[2]  & ((~new_n460_ ^ \a[5] ) ^ ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] ))))) | ((~\a[2]  | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )) | (new_n462_ & (~new_n461_ ^ \a[5] ))) & (new_n531_ | (\a[2]  & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )) & (~new_n462_ | (new_n461_ ^ \a[5] ))) | (~\a[2]  & (new_n462_ ^ (new_n461_ ^ \a[5] ))))))))) | (\a[2]  & ((new_n458_ & \a[5] ) | (~new_n458_ & ~\a[5] ) | ((~new_n459_ | ~\a[5] ) & ((new_n459_ & \a[5] ) | (~new_n459_ & ~\a[5] ) | ((~new_n460_ | ~\a[5] ) & ((new_n460_ & \a[5] ) | (~new_n460_ & ~\a[5] ) | ((~new_n461_ | ~\a[5] ) & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )))))))) & ((new_n458_ ^ \a[5] ) | (new_n459_ & \a[5] ) | ((~new_n459_ | ~\a[5] ) & (new_n459_ | \a[5] ) & ((new_n460_ & \a[5] ) | ((~new_n460_ | ~\a[5] ) & (new_n460_ | \a[5] ) & ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )))))))) | (~\a[2]  & ((~new_n458_ ^ \a[5] ) ^ ((new_n459_ & \a[5] ) | ((~new_n459_ | ~\a[5] ) & (new_n459_ | \a[5] ) & ((new_n460_ & \a[5] ) | ((~new_n460_ | ~\a[5] ) & (new_n460_ | \a[5] ) & ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] ))))))))));
  assign new_n531_ = (~new_n532_ | ~\a[2] ) & ((~new_n532_ & ~\a[2] ) | (new_n532_ & \a[2] ) | ((~\a[2]  | (new_n587_ & (new_n585_ | (~new_n464_ & new_n586_))) | (~new_n587_ & ~new_n585_ & (new_n464_ | ~new_n586_))) & (((~\a[2]  | (new_n464_ & ~new_n586_) | (~new_n464_ & new_n586_)) & (new_n533_ | (\a[2]  & (~new_n464_ | new_n586_) & (new_n464_ | ~new_n586_)) | (~\a[2]  & (~new_n464_ ^ ~new_n586_)))) | (\a[2]  & (~new_n587_ | (~new_n585_ & (new_n464_ | ~new_n586_))) & (new_n587_ | new_n585_ | (~new_n464_ & new_n586_))) | (~\a[2]  & (~new_n587_ ^ (new_n585_ | (~new_n464_ & new_n586_)))))));
  assign new_n532_ = (~new_n463_ ^ ~\a[5] ) ^ ((\a[5]  & ((new_n324_ & \a[8] ) | (~new_n324_ & ~\a[8] ) | ((~new_n325_ | ~\a[8] ) & ((new_n325_ & \a[8] ) | (~new_n325_ & ~\a[8] ) | ((~new_n326_ | ~\a[8] ) & (new_n328_ | (new_n326_ & \a[8] ) | (~new_n326_ & ~\a[8] )))))) & ((new_n324_ ^ \a[8] ) | (new_n325_ & \a[8] ) | ((~new_n325_ | ~\a[8] ) & (new_n325_ | \a[8] ) & ((new_n326_ & \a[8] ) | (~new_n328_ & (~new_n326_ | ~\a[8] ) & (new_n326_ | \a[8] )))))) | ((~\a[5]  | ((~new_n324_ | ~\a[8] ) & (new_n324_ | \a[8] ) & ((new_n325_ & \a[8] ) | ((~new_n325_ | ~\a[8] ) & (new_n325_ | \a[8] ) & ((new_n326_ & \a[8] ) | (~new_n328_ & (~new_n326_ | ~\a[8] ) & (new_n326_ | \a[8] )))))) | ((~new_n324_ ^ \a[8] ) & (~new_n325_ | ~\a[8] ) & ((new_n325_ & \a[8] ) | (~new_n325_ & ~\a[8] ) | ((~new_n326_ | ~\a[8] ) & (new_n328_ | (new_n326_ & \a[8] ) | (~new_n326_ & ~\a[8] )))))) & (\a[5]  | ((new_n324_ ^ \a[8] ) ^ ((new_n325_ & \a[8] ) | ((~new_n325_ | ~\a[8] ) & (new_n325_ | \a[8] ) & ((new_n326_ & \a[8] ) | (~new_n328_ & (~new_n326_ | ~\a[8] ) & (new_n326_ | \a[8] ))))))) & ((\a[5]  & ((new_n325_ & \a[8] ) | (~new_n325_ & ~\a[8] ) | ((~new_n326_ | ~\a[8] ) & (new_n328_ | (new_n326_ & \a[8] ) | (~new_n326_ & ~\a[8] )))) & ((new_n325_ ^ \a[8] ) | (new_n326_ & \a[8] ) | (~new_n328_ & (~new_n326_ | ~\a[8] ) & (new_n326_ | \a[8] )))) | (~new_n464_ & (~\a[5]  | ((~new_n325_ | ~\a[8] ) & (new_n325_ | \a[8] ) & ((new_n326_ & \a[8] ) | (~new_n328_ & (~new_n326_ | ~\a[8] ) & (new_n326_ | \a[8] )))) | ((~new_n325_ ^ \a[8] ) & (~new_n326_ | ~\a[8] ) & (new_n328_ | (new_n326_ & \a[8] ) | (~new_n326_ & ~\a[8] )))) & (\a[5]  | ((new_n325_ ^ \a[8] ) ^ ((new_n326_ & \a[8] ) | (~new_n328_ & (~new_n326_ | ~\a[8] ) & (new_n326_ | \a[8] )))))))));
  assign new_n533_ = (~new_n534_ | ~\a[2] ) & ((~new_n534_ & ~\a[2] ) | (new_n534_ & \a[2] ) | ((~\a[2]  | ((~new_n466_ | ~\a[5] ) & (new_n466_ | \a[5] ) & ((new_n467_ & \a[5] ) | ((~new_n467_ | ~\a[5] ) & (new_n467_ | \a[5] ) & ((new_n468_ & \a[5] ) | (~new_n470_ & (~new_n468_ | ~\a[5] ) & (new_n468_ | \a[5] )))))) | ((~new_n466_ ^ \a[5] ) & (~new_n467_ | ~\a[5] ) & ((new_n467_ & \a[5] ) | (~new_n467_ & ~\a[5] ) | ((~new_n468_ | ~\a[5] ) & (new_n470_ | (new_n468_ & \a[5] ) | (~new_n468_ & ~\a[5] )))))) & ((\a[2]  & ((new_n466_ & \a[5] ) | (~new_n466_ & ~\a[5] ) | ((~new_n467_ | ~\a[5] ) & ((new_n467_ & \a[5] ) | (~new_n467_ & ~\a[5] ) | ((~new_n468_ | ~\a[5] ) & (new_n470_ | (new_n468_ & \a[5] ) | (~new_n468_ & ~\a[5] )))))) & ((new_n466_ ^ \a[5] ) | (new_n467_ & \a[5] ) | ((~new_n467_ | ~\a[5] ) & (new_n467_ | \a[5] ) & ((new_n468_ & \a[5] ) | (~new_n470_ & (~new_n468_ | ~\a[5] ) & (new_n468_ | \a[5] )))))) | (~\a[2]  & ((~new_n466_ ^ \a[5] ) ^ ((new_n467_ & \a[5] ) | ((~new_n467_ | ~\a[5] ) & (new_n467_ | \a[5] ) & ((new_n468_ & \a[5] ) | (~new_n470_ & (~new_n468_ | ~\a[5] ) & (new_n468_ | \a[5] ))))))) | ((~\a[2]  | ((~new_n467_ | ~\a[5] ) & (new_n467_ | \a[5] ) & ((new_n468_ & \a[5] ) | (~new_n470_ & (~new_n468_ | ~\a[5] ) & (new_n468_ | \a[5] )))) | ((~new_n467_ ^ \a[5] ) & (~new_n468_ | ~\a[5] ) & (new_n470_ | (new_n468_ & \a[5] ) | (~new_n468_ & ~\a[5] )))) & (new_n535_ | (\a[2]  & ((new_n467_ & \a[5] ) | (~new_n467_ & ~\a[5] ) | ((~new_n468_ | ~\a[5] ) & (new_n470_ | (new_n468_ & \a[5] ) | (~new_n468_ & ~\a[5] )))) & ((new_n467_ ^ \a[5] ) | (new_n468_ & \a[5] ) | (~new_n470_ & (~new_n468_ | ~\a[5] ) & (new_n468_ | \a[5] )))) | (~\a[2]  & ((~new_n467_ ^ \a[5] ) ^ ((new_n468_ & \a[5] ) | (~new_n470_ & (~new_n468_ | ~\a[5] ) & (new_n468_ | \a[5] ))))))))));
  assign new_n534_ = ((new_n466_ & \a[5] ) | ((~new_n466_ | ~\a[5] ) & (new_n466_ | \a[5] ) & ((new_n467_ & \a[5] ) | (((new_n468_ & \a[5] ) | (~new_n470_ & (new_n468_ | \a[5] ) & (~new_n468_ | ~\a[5] ))) & (~new_n467_ | ~\a[5] ) & (new_n467_ | \a[5] ))))) ^ (\a[5]  ^ (new_n328_ ^ ~new_n465_));
  assign new_n535_ = (~\a[2]  | (new_n583_ & ~new_n537_ & ~new_n538_)) & ((new_n470_ & ~new_n536_) | (~new_n470_ & new_n536_) | (~\a[2]  & (~new_n537_ | ~new_n538_ | ~new_n584_)));
  assign new_n536_ = \a[5]  ^ (new_n469_ ^ ~new_n331_);
  assign new_n537_ = (new_n472_ ^ \a[5] ) ^ ((\a[5]  & (((~new_n334_ | ~\a[8] ) & ((new_n334_ & \a[8] ) | (~new_n334_ & ~\a[8] ) | ((~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] ))))) | (new_n471_ & \a[8] ) | (~new_n471_ & ~\a[8] )) & ((new_n334_ & \a[8] ) | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))) | (new_n471_ ^ \a[8] ))) | ((~\a[5]  | (((new_n334_ & \a[8] ) | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] ))))) & (~new_n471_ | ~\a[8] ) & (new_n471_ | \a[8] )) | ((~new_n334_ | ~\a[8] ) & ((new_n334_ & \a[8] ) | (~new_n334_ & ~\a[8] ) | ((~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))) & (~new_n471_ ^ \a[8] ))) & (\a[5]  | (((new_n334_ & \a[8] ) | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] ))))) ^ (new_n471_ ^ \a[8] ))) & ((\a[5]  & ((new_n334_ & \a[8] ) | (~new_n334_ & ~\a[8] ) | ((~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))) & ((new_n334_ ^ \a[8] ) | (new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))) | (~new_n473_ & (~\a[5]  | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))) | ((~new_n334_ ^ \a[8] ) & (~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))) & (\a[5]  | ((new_n334_ ^ \a[8] ) ^ ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))))))));
  assign new_n538_ = (new_n582_ ^ \a[2] ) & ((new_n539_ & \a[2] ) | (~new_n540_ & (new_n539_ | \a[2] ) & (~new_n539_ | ~\a[2] )));
  assign new_n539_ = (new_n475_ ^ \a[5] ) ^ ((new_n477_ & \a[5] ) | (((new_n478_ & \a[5] ) | (~new_n480_ & (new_n478_ | \a[5] ) & (~new_n478_ | ~\a[5] ))) & (~new_n477_ | ~\a[5] ) & (new_n477_ | \a[5] )));
  assign new_n540_ = (~\a[2]  | ((~new_n477_ | ~\a[5] ) & (new_n477_ | \a[5] ) & ((new_n478_ & \a[5] ) | (~new_n480_ & (~new_n478_ | ~\a[5] ) & (new_n478_ | \a[5] )))) | ((~new_n477_ ^ \a[5] ) & (~new_n478_ | ~\a[5] ) & (new_n480_ | (new_n478_ & \a[5] ) | (~new_n478_ & ~\a[5] )))) & (((~\a[2]  | (~new_n480_ & (~new_n478_ | ~\a[5] ) & (new_n478_ | \a[5] )) | (new_n480_ & (~new_n478_ ^ \a[5] ))) & (((~new_n541_ | ~\a[2] ) & (((~new_n543_ | ~\a[2] ) & (new_n544_ | (~new_n543_ & ~\a[2] ) | (new_n543_ & \a[2] ))) | (new_n541_ & \a[2] ) | (~new_n541_ & ~\a[2] ))) | (\a[2]  & (new_n480_ | (new_n478_ & \a[5] ) | (~new_n478_ & ~\a[5] )) & (~new_n480_ | (new_n478_ ^ \a[5] ))) | (~\a[2]  & (new_n480_ ^ (new_n478_ ^ \a[5] ))))) | (\a[2]  & ((new_n477_ & \a[5] ) | (~new_n477_ & ~\a[5] ) | ((~new_n478_ | ~\a[5] ) & (new_n480_ | (new_n478_ & \a[5] ) | (~new_n478_ & ~\a[5] )))) & ((new_n477_ ^ \a[5] ) | (new_n478_ & \a[5] ) | (~new_n480_ & (~new_n478_ | ~\a[5] ) & (new_n478_ | \a[5] )))) | (~\a[2]  & ((~new_n477_ ^ \a[5] ) ^ ((new_n478_ & \a[5] ) | (~new_n480_ & (~new_n478_ | ~\a[5] ) & (new_n478_ | \a[5] ))))));
  assign new_n541_ = new_n542_ ^ (new_n482_ | (~new_n482_ & ~new_n519_ & ((~new_n521_ & (new_n349_ | ~new_n372_) & (~new_n349_ | new_n372_)) | (~new_n484_ & (new_n521_ | (~new_n349_ & new_n372_) | (new_n349_ & ~new_n372_)) & (~new_n521_ | (~new_n349_ ^ new_n372_))))));
  assign new_n542_ = ~new_n520_ ^ ((new_n344_ | (new_n373_ & (new_n346_ | (~new_n349_ & new_n372_)))) ^ (new_n342_ ^ ~new_n374_));
  assign new_n543_ = (~new_n482_ & ~new_n519_) ^ ((~new_n521_ & (~new_n349_ | new_n372_) & (new_n349_ | ~new_n372_)) | (~new_n484_ & (~new_n521_ | (new_n349_ ^ ~new_n372_)) & (new_n521_ | (new_n349_ & ~new_n372_) | (~new_n349_ & new_n372_))));
  assign new_n544_ = (~\a[2]  | (new_n484_ & ~new_n545_) | (~new_n484_ & new_n545_)) & ((\a[2]  & (~new_n484_ | new_n545_) & (new_n484_ | ~new_n545_)) | (~\a[2]  & (~new_n484_ ^ ~new_n545_)) | ((~new_n546_ | new_n581_) & ((new_n546_ & ~new_n581_) | (~new_n546_ & new_n581_) | (~new_n547_ & (new_n549_ | ~new_n580_)))));
  assign new_n545_ = ~new_n521_ ^ (new_n349_ ^ ~new_n372_);
  assign new_n546_ = (new_n487_ | (new_n517_ & (new_n489_ | (~new_n492_ & new_n516_)))) ^ (new_n485_ ^ ~new_n518_);
  assign new_n547_ = ~new_n548_ & (~new_n517_ | (~new_n489_ & (new_n492_ | ~new_n516_))) & (new_n517_ | new_n489_ | (~new_n492_ & new_n516_));
  assign new_n548_ = \a[2]  ^ (((~\b[14]  ^ ((\b[13]  & \b[14] ) | (~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[14]  | \a[0]  | ~\a[1] ) & (~\b[13]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ));
  assign new_n549_ = (new_n578_ | (new_n492_ & ~new_n516_) | (~new_n492_ & new_n516_)) & (((~new_n550_ | new_n579_) & ((~new_n552_ & (new_n554_ | ~new_n577_)) | (new_n550_ & ~new_n579_) | (~new_n550_ & new_n579_))) | (~new_n578_ & (~new_n492_ | new_n516_) & (new_n492_ | ~new_n516_)) | (new_n578_ & (~new_n492_ ^ ~new_n516_)));
  assign new_n550_ = new_n551_ ^ (new_n495_ | (new_n497_ & ((~new_n515_ & (new_n360_ | (~new_n359_ & new_n367_) | (new_n359_ & ~new_n367_)) & (~new_n360_ | (~new_n359_ ^ new_n367_))) | (~new_n498_ & (new_n515_ | (~new_n360_ & (new_n359_ | ~new_n367_) & (~new_n359_ | new_n367_)) | (new_n360_ & (new_n359_ ^ new_n367_))) & (~new_n515_ | (~new_n360_ ^ (~new_n359_ ^ new_n367_)))))));
  assign new_n551_ = ~new_n513_ ^ ((new_n355_ ^ ~new_n356_) ^ ((new_n357_ & ~new_n358_) | ((new_n357_ | ~new_n358_) & (~new_n357_ | new_n358_) & ((~new_n359_ & new_n367_) | (~new_n360_ & (new_n359_ | ~new_n367_) & (~new_n359_ | new_n367_))))));
  assign new_n552_ = ~new_n553_ & (~new_n497_ | ((new_n515_ | (~new_n360_ & (new_n359_ | ~new_n367_) & (~new_n359_ | new_n367_)) | (new_n360_ & (new_n359_ ^ new_n367_))) & (new_n498_ | (~new_n515_ & (new_n360_ | (~new_n359_ & new_n367_) | (new_n359_ & ~new_n367_)) & (~new_n360_ | (~new_n359_ ^ new_n367_))) | (new_n515_ & (new_n360_ ^ (~new_n359_ ^ new_n367_)))))) & (new_n497_ | (~new_n515_ & (new_n360_ | (~new_n359_ & new_n367_) | (new_n359_ & ~new_n367_)) & (~new_n360_ | (~new_n359_ ^ new_n367_))) | (~new_n498_ & (new_n515_ | (~new_n360_ & (new_n359_ | ~new_n367_) & (~new_n359_ | new_n367_)) | (new_n360_ & (new_n359_ ^ new_n367_))) & (~new_n515_ | (~new_n360_ ^ (~new_n359_ ^ new_n367_)))));
  assign new_n553_ = \a[2]  ^ ((~new_n106_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[10]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[11]  | \a[0]  | ~\a[1] ) & (~\b[12]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )));
  assign new_n554_ = (new_n556_ | (new_n498_ & ~new_n555_) | (~new_n498_ & new_n555_)) & ((~new_n556_ & (~new_n498_ | new_n555_) & (new_n498_ | ~new_n555_)) | (new_n556_ & (~new_n498_ ^ ~new_n555_)) | ((~new_n557_ | new_n576_) & ((~new_n558_ & (new_n560_ | ~new_n575_)) | (new_n557_ & ~new_n576_) | (~new_n557_ & new_n576_))));
  assign new_n555_ = ~new_n515_ ^ (~new_n360_ ^ (new_n359_ ^ ~new_n367_));
  assign new_n556_ = \a[2]  ^ ((~new_n112_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[9]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[10]  | \a[0]  | ~\a[1] ) & (~\b[11]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )));
  assign new_n557_ = (new_n499_ ^ ~new_n500_) ^ ((new_n501_ & ~new_n502_) | ((new_n501_ | ~new_n502_) & (~new_n501_ | new_n502_) & ((~new_n503_ & new_n512_) | (~new_n506_ & (new_n503_ | ~new_n512_) & (~new_n503_ | new_n512_)))));
  assign new_n558_ = ~new_n559_ & ((new_n501_ & ~new_n502_) | (~new_n501_ & new_n502_) | ((new_n503_ | ~new_n512_) & (new_n506_ | (~new_n503_ & new_n512_) | (new_n503_ & ~new_n512_)))) & ((new_n501_ ^ ~new_n502_) | (~new_n503_ & new_n512_) | (~new_n506_ & (new_n503_ | ~new_n512_) & (~new_n503_ | new_n512_)));
  assign new_n559_ = \a[2]  ^ ((~\b[7]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[8]  | \a[0]  | ~\a[1] ) & (~\b[9]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))));
  assign new_n560_ = (new_n562_ | (new_n506_ & ~new_n561_) | (~new_n506_ & new_n561_)) & ((~new_n562_ & (~new_n506_ | new_n561_) & (new_n506_ | ~new_n561_)) | (new_n562_ & (~new_n506_ ^ ~new_n561_)) | ((new_n563_ | ~new_n564_) & ((new_n563_ & ~new_n564_) | (~new_n563_ & new_n564_) | ((new_n565_ | ~new_n568_) & (new_n569_ | (~new_n565_ & new_n568_) | (new_n565_ & ~new_n568_))))));
  assign new_n561_ = new_n512_ ^ (~\a[5]  ^ (new_n505_ & (~new_n63_ | ~new_n504_)));
  assign new_n562_ = \a[2]  ^ ((~\b[6]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[7]  | \a[0]  | ~\a[1] ) & (~\b[8]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n80_ & (~\b[7]  ^ \b[8] ))));
  assign new_n563_ = \a[2]  ^ ((~new_n75_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[5]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[6]  | \a[0]  | ~\a[1] ) & (~\b[7]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )));
  assign new_n564_ = (new_n509_ | (~new_n510_ & new_n511_)) ^ (new_n508_ ^ (~\a[5]  ^ (new_n507_ & (~new_n66_ | ~new_n504_))));
  assign new_n565_ = \a[2]  ^ (new_n567_ & (~new_n60_ | ~new_n566_));
  assign new_n566_ = \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] );
  assign new_n567_ = (~\b[4]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[6]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[5]  | \a[0]  | ~\a[1] );
  assign new_n568_ = new_n510_ ^ ~new_n511_;
  assign new_n569_ = (~new_n571_ | (\a[2]  ^ (new_n570_ & (~new_n63_ | ~new_n566_)))) & ((new_n571_ & (~\a[2]  ^ (new_n570_ & (~new_n63_ | ~new_n566_)))) | (~new_n571_ & (~\a[2]  | ~new_n570_ | (new_n63_ & new_n566_)) & (\a[2]  | (new_n570_ & (~new_n63_ | ~new_n566_)))) | ((new_n572_ | ~new_n573_) & (new_n574_ | (~new_n572_ & new_n573_) | (new_n572_ & ~new_n573_))));
  assign new_n570_ = (~\b[3]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[5]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[4]  | \a[0]  | ~\a[1] );
  assign new_n571_ = (~\a[5]  | ((~\b[0]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )))) ^ ((~\b[1]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[2]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )));
  assign new_n572_ = \a[2]  ^ ((~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )))) | ((~\b[3]  ^ \b[4] ) & (~\b[2]  | ~\b[3] ) & ((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[4]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[3]  | \a[0]  | ~\a[1] ));
  assign new_n573_ = ((\b[0]  & (\a[2]  ^ ~\a[3] ) & (\a[3]  | \a[4] ) & (~\a[3]  | ~\a[4] )) | (\b[1]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (\a[4]  ^ ~\a[5] )) | ((\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (\a[4]  | \a[5] ) & (~\a[4]  | ~\a[5] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[5]  & \b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ));
  assign new_n574_ = (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[2]  ^ ((~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] ) & (((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))))) & (((~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\a[2]  | (\b[1]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[3]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[2]  & ~\a[0]  & \a[1] ) | (((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )) & ((\b[2]  ^ \b[3] ) | (\b[1]  & (\b[0]  | \b[2] ))) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] ))) & (\a[2]  | ((~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] ) & (((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))))) | ~\a[2]  | (\b[1]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[0]  & ~\a[0]  & \a[1] ) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\a[0]  & \b[0] ) | (\b[2]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[1]  & ~\a[0]  & \a[1] ) | (\b[0]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | ((~\b[2]  ^ (\b[0]  | ~\b[1] )) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )));
  assign new_n575_ = ~new_n559_ ^ ((new_n501_ ^ ~new_n502_) ^ ((~new_n503_ & new_n512_) | (~new_n506_ & (new_n503_ | ~new_n512_) & (~new_n503_ | new_n512_))));
  assign new_n576_ = \a[2]  ^ ((((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n80_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n80_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[8]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[10]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[9]  | \a[0]  | ~\a[1] ));
  assign new_n577_ = ~new_n553_ ^ (new_n497_ ^ ((~new_n515_ & (new_n360_ | (~new_n359_ & new_n367_) | (new_n359_ & ~new_n367_)) & (~new_n360_ | (~new_n359_ ^ new_n367_))) | (~new_n498_ & (new_n515_ | (~new_n360_ & (new_n359_ | ~new_n367_) & (~new_n359_ | new_n367_)) | (new_n360_ & (new_n359_ ^ new_n367_))) & (~new_n515_ | (~new_n360_ ^ (~new_n359_ ^ new_n367_))))));
  assign new_n578_ = \a[2]  ^ ((~\b[12]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[13]  | \a[0]  | ~\a[1] ) & (~\b[14]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | (~new_n114_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n114_ & (~\b[13]  ^ \b[14] ))));
  assign new_n579_ = \a[2]  ^ ((~new_n149_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[11]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[12]  | \a[0]  | ~\a[1] ) & (~\b[13]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )));
  assign new_n580_ = ~new_n548_ ^ (new_n517_ ^ (new_n489_ | (~new_n492_ & new_n516_)));
  assign new_n581_ = \a[2]  ^ (~\b[14]  | (((~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (new_n164_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))));
  assign new_n582_ = ((new_n475_ & \a[5] ) | ((~new_n475_ | ~\a[5] ) & (new_n475_ | \a[5] ) & ((new_n477_ & \a[5] ) | (((new_n478_ & \a[5] ) | (~new_n480_ & (new_n478_ | \a[5] ) & (~new_n478_ | ~\a[5] ))) & (~new_n477_ | ~\a[5] ) & (new_n477_ | \a[5] ))))) ^ (\a[5]  ^ (new_n337_ ^ ~new_n474_));
  assign new_n583_ = (((~\a[5]  | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))) | ((~new_n334_ ^ \a[8] ) & (~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))) & (new_n473_ | (\a[5]  & ((new_n334_ & \a[8] ) | (~new_n334_ & ~\a[8] ) | ((~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))) & ((new_n334_ ^ \a[8] ) | (new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))) | (~\a[5]  & ((~new_n334_ ^ \a[8] ) ^ ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] ))))))) ^ (\a[5]  ^ (((new_n334_ & \a[8] ) | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] ))))) ^ (new_n471_ ^ \a[8] )))) & ~new_n582_ & (new_n473_ ^ (\a[5]  ^ ((new_n334_ ^ \a[8] ) ^ ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] ))))));
  assign new_n584_ = ((\a[5]  & ((~new_n471_ & ~\a[8] ) | (new_n471_ & \a[8] ) | ((~new_n334_ | ~\a[8] ) & ((new_n334_ & \a[8] ) | (~new_n334_ & ~\a[8] ) | ((~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))))) & ((~new_n471_ ^ ~\a[8] ) | (new_n334_ & \a[8] ) | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))))) | (~\a[5]  & ((new_n471_ ^ ~\a[8] ) ^ ((new_n334_ & \a[8] ) | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] ))))))) | ((~\a[5]  | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))) | ((~new_n334_ ^ \a[8] ) & (~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))) & (new_n473_ | (\a[5]  & ((new_n334_ & \a[8] ) | (~new_n334_ & ~\a[8] ) | ((~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))) & ((new_n334_ ^ \a[8] ) | (new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))) | (~\a[5]  & ((~new_n334_ ^ \a[8] ) ^ ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))))))) & ((\a[5]  ^ ((~new_n471_ ^ ~\a[8] ) ^ ((new_n334_ & \a[8] ) | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] ))))))) | (\a[5]  & ((new_n334_ & \a[8] ) | (~new_n334_ & ~\a[8] ) | ((~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))) & ((new_n334_ ^ \a[8] ) | (new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))) | (~new_n473_ & (~\a[5]  | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))) | ((~new_n334_ ^ \a[8] ) & (~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))) & (\a[5]  | ((new_n334_ ^ \a[8] ) ^ ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] ))))))) & (new_n473_ | (\a[5]  & ((new_n334_ & \a[8] ) | (~new_n334_ & ~\a[8] ) | ((~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))) & ((new_n334_ ^ \a[8] ) | (new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))) | (~\a[5]  & ((~new_n334_ ^ \a[8] ) ^ ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))))) & (~new_n473_ | (\a[5]  ^ ((new_n334_ ^ \a[8] ) ^ ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] ))))));
  assign new_n585_ = \a[5]  & ((new_n325_ & \a[8] ) | (~new_n325_ & ~\a[8] ) | ((~new_n326_ | ~\a[8] ) & (new_n328_ | (new_n326_ & \a[8] ) | (~new_n326_ & ~\a[8] )))) & ((new_n325_ ^ \a[8] ) | (new_n326_ & \a[8] ) | (~new_n328_ & (~new_n326_ | ~\a[8] ) & (new_n326_ | \a[8] )));
  assign new_n586_ = \a[5]  ^ ((new_n325_ ^ \a[8] ) ^ ((new_n326_ & \a[8] ) | (~new_n328_ & (~new_n326_ | ~\a[8] ) & (new_n326_ | \a[8] ))));
  assign new_n587_ = \a[5]  ^ ((new_n324_ ^ \a[8] ) ^ ((new_n325_ & \a[8] ) | ((~new_n325_ | ~\a[8] ) & (new_n325_ | \a[8] ) & ((new_n326_ & \a[8] ) | (~new_n328_ & (~new_n326_ | ~\a[8] ) & (new_n326_ | \a[8] ))))));
  assign new_n588_ = (\a[5]  ^ (new_n453_ ^ ~new_n457_)) ^ ((new_n458_ & \a[5] ) | ((~new_n458_ | ~\a[5] ) & (new_n458_ | \a[5] ) & ((new_n459_ & \a[5] ) | ((~new_n459_ | ~\a[5] ) & (new_n459_ | \a[5] ) & ((new_n460_ & \a[5] ) | ((~new_n460_ | ~\a[5] ) & (new_n460_ | \a[5] ) & ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )))))))));
  assign new_n589_ = ((~\a[2]  ^ (new_n526_ ^ ~new_n528_)) ^ ((new_n529_ & \a[2] ) | ((~new_n529_ | ~\a[2] ) & (new_n529_ | \a[2] ) & ((new_n588_ & \a[2] ) | (~new_n530_ & (~new_n588_ | ~\a[2] ) & (new_n588_ | \a[2] )))))) & ((~new_n529_ ^ \a[2] ) ^ ((new_n588_ & \a[2] ) | (~new_n530_ & (~new_n588_ | ~\a[2] ) & (new_n588_ | \a[2] )))) & ~new_n590_ & new_n591_ & (new_n530_ ^ (new_n588_ ^ \a[2] ));
  assign new_n590_ = ((\a[2]  & ((new_n459_ & \a[5] ) | (~new_n459_ & ~\a[5] ) | ((~new_n460_ | ~\a[5] ) & ((new_n460_ & \a[5] ) | (~new_n460_ & ~\a[5] ) | ((~new_n461_ | ~\a[5] ) & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )))))) & ((new_n459_ ^ \a[5] ) | (new_n460_ & \a[5] ) | ((~new_n460_ | ~\a[5] ) & (new_n460_ | \a[5] ) & ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )))))) | ((~\a[2]  | ((~new_n459_ | ~\a[5] ) & (new_n459_ | \a[5] ) & ((new_n460_ & \a[5] ) | ((~new_n460_ | ~\a[5] ) & (new_n460_ | \a[5] ) & ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )))))) | ((~new_n459_ ^ \a[5] ) & (~new_n460_ | ~\a[5] ) & ((new_n460_ & \a[5] ) | (~new_n460_ & ~\a[5] ) | ((~new_n461_ | ~\a[5] ) & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )))))) & (\a[2]  | ((new_n459_ ^ \a[5] ) ^ ((new_n460_ & \a[5] ) | ((~new_n460_ | ~\a[5] ) & (new_n460_ | \a[5] ) & ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] ))))))) & ((\a[2]  & ((new_n460_ & \a[5] ) | (~new_n460_ & ~\a[5] ) | ((~new_n461_ | ~\a[5] ) & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )))) & ((new_n460_ ^ \a[5] ) | (new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )))) | ((~\a[2]  | ((~new_n460_ | ~\a[5] ) & (new_n460_ | \a[5] ) & ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )))) | ((~new_n460_ ^ \a[5] ) & (~new_n461_ | ~\a[5] ) & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )))) & (\a[2]  | ((new_n460_ ^ \a[5] ) ^ ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] ))))) & ((\a[2]  & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )) & (~new_n462_ | (new_n461_ ^ \a[5] ))) | (~new_n531_ & (~\a[2]  | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )) | (new_n462_ & (~new_n461_ ^ \a[5] ))) & (\a[2]  | (~new_n462_ ^ (new_n461_ ^ \a[5] ))))))))) ^ (\a[2]  ^ ((new_n458_ ^ \a[5] ) ^ ((new_n459_ & \a[5] ) | ((~new_n459_ | ~\a[5] ) & (new_n459_ | \a[5] ) & ((new_n460_ & \a[5] ) | ((~new_n460_ | ~\a[5] ) & (new_n460_ | \a[5] ) & ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )))))))));
  assign new_n591_ = ((~\a[2]  ^ ((new_n459_ ^ \a[5] ) ^ ((new_n460_ & \a[5] ) | ((~new_n460_ | ~\a[5] ) & (new_n460_ | \a[5] ) & ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] ))))))) ^ ((\a[2]  & ((new_n460_ & \a[5] ) | (~new_n460_ & ~\a[5] ) | ((~new_n461_ | ~\a[5] ) & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )))) & ((new_n460_ ^ \a[5] ) | (new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )))) | ((~\a[2]  | ((~new_n460_ | ~\a[5] ) & (new_n460_ | \a[5] ) & ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )))) | ((~new_n460_ ^ \a[5] ) & (~new_n461_ | ~\a[5] ) & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )))) & (\a[2]  | ((new_n460_ ^ \a[5] ) ^ ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] ))))) & ((\a[2]  & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )) & (~new_n462_ | (new_n461_ ^ \a[5] ))) | (~new_n531_ & (~\a[2]  | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )) | (new_n462_ & (~new_n461_ ^ \a[5] ))) & (\a[2]  | (~new_n462_ ^ (new_n461_ ^ \a[5] )))))))) & ((~\a[2]  ^ ((new_n460_ ^ \a[5] ) ^ ((new_n461_ & \a[5] ) | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] ))))) ^ ((\a[2]  & (new_n462_ | (new_n461_ & \a[5] ) | (~new_n461_ & ~\a[5] )) & (~new_n462_ | (new_n461_ ^ \a[5] ))) | (~new_n531_ & (~\a[2]  | (~new_n462_ & (~new_n461_ | ~\a[5] ) & (new_n461_ | \a[5] )) | (new_n462_ & (~new_n461_ ^ \a[5] ))) & (\a[2]  | (~new_n462_ ^ (new_n461_ ^ \a[5] )))))) & new_n592_ & (new_n531_ ^ (\a[2]  ^ (~new_n462_ ^ (new_n461_ ^ \a[5] ))));
  assign new_n592_ = ((~new_n532_ ^ \a[2] ) ^ ((\a[2]  & (~new_n587_ | (~new_n585_ & (new_n464_ | ~new_n586_))) & (new_n587_ | new_n585_ | (~new_n464_ & new_n586_))) | (((\a[2]  & (new_n464_ | ~new_n586_) & (~new_n464_ | new_n586_)) | (~new_n533_ & (~\a[2]  | (~new_n464_ & new_n586_) | (new_n464_ & ~new_n586_)) & (\a[2]  | (~new_n464_ ^ new_n586_)))) & (~\a[2]  | (new_n587_ & (new_n585_ | (~new_n464_ & new_n586_))) | (~new_n587_ & ~new_n585_ & (new_n464_ | ~new_n586_))) & (\a[2]  | (new_n587_ ^ (new_n585_ | (~new_n464_ & new_n586_))))))) & (((~\a[2]  | (~new_n464_ & new_n586_) | (new_n464_ & ~new_n586_)) & (new_n533_ | (\a[2]  & (new_n464_ | ~new_n586_) & (~new_n464_ | new_n586_)) | (~\a[2]  & (new_n464_ ^ new_n586_)))) ^ (\a[2]  ^ (new_n587_ ^ (new_n585_ | (~new_n464_ & new_n586_))))) & new_n593_ & (new_n533_ ^ (\a[2]  ^ (~new_n464_ ^ new_n586_)));
  assign new_n593_ = (~new_n599_ ^ (new_n594_ | (~new_n594_ & ~new_n598_ & (new_n595_ | (~new_n535_ & ~new_n595_ & ~new_n596_))))) & ((new_n594_ | new_n598_) ^ (new_n595_ | (~new_n535_ & ~new_n595_ & ~new_n596_))) & (~new_n535_ | (~new_n595_ & ~new_n596_)) & new_n597_ & new_n600_ & (new_n535_ | new_n595_ | new_n596_);
  assign new_n594_ = \a[2]  & ((new_n466_ & \a[5] ) | (~new_n466_ & ~\a[5] ) | ((~new_n467_ | ~\a[5] ) & ((new_n467_ & \a[5] ) | (~new_n467_ & ~\a[5] ) | ((~new_n468_ | ~\a[5] ) & (new_n470_ | (new_n468_ & \a[5] ) | (~new_n468_ & ~\a[5] )))))) & ((new_n466_ ^ \a[5] ) | (new_n467_ & \a[5] ) | ((~new_n467_ | ~\a[5] ) & (new_n467_ | \a[5] ) & ((new_n468_ & \a[5] ) | (~new_n470_ & (~new_n468_ | ~\a[5] ) & (new_n468_ | \a[5] )))));
  assign new_n595_ = \a[2]  & ((new_n467_ & \a[5] ) | (~new_n467_ & ~\a[5] ) | ((~new_n468_ | ~\a[5] ) & (new_n470_ | (new_n468_ & \a[5] ) | (~new_n468_ & ~\a[5] )))) & ((new_n467_ ^ \a[5] ) | (new_n468_ & \a[5] ) | (~new_n470_ & (~new_n468_ | ~\a[5] ) & (new_n468_ | \a[5] )));
  assign new_n596_ = ~\a[2]  & ((~new_n467_ ^ \a[5] ) ^ ((new_n468_ & \a[5] ) | (~new_n470_ & new_n536_)));
  assign new_n597_ = new_n470_ ^ ~new_n536_;
  assign new_n598_ = ~\a[2]  & ((new_n466_ ^ ~\a[5] ) ^ ((new_n467_ & \a[5] ) | ((~new_n467_ | ~\a[5] ) & (new_n467_ | \a[5] ) & ((new_n468_ & \a[5] ) | (~new_n470_ & new_n536_)))));
  assign new_n599_ = \a[2]  ^ (((new_n466_ & \a[5] ) | ((~new_n466_ | ~\a[5] ) & (new_n466_ | \a[5] ) & ((new_n467_ & \a[5] ) | ((~new_n467_ | ~\a[5] ) & (new_n467_ | \a[5] ) & ((new_n468_ & \a[5] ) | (~new_n470_ & (~new_n468_ | ~\a[5] ) & (new_n468_ | \a[5] ))))))) ^ (\a[5]  ^ (new_n328_ ^ ~new_n465_)));
  assign new_n600_ = ~new_n537_ & ((~new_n582_ ^ \a[2] ) | ((~new_n539_ | ~\a[2] ) & (new_n540_ | (new_n539_ & \a[2] ) | (~new_n539_ & ~\a[2] )))) & ((~new_n582_ & \a[2] ) | (new_n582_ & ~\a[2] ) | (new_n539_ & \a[2] ) | (~new_n540_ & (~new_n539_ | ~\a[2] ) & (new_n539_ | \a[2] ))) & new_n602_ & new_n601_ & (new_n540_ ^ (new_n539_ ^ \a[2] ));
  assign new_n601_ = (\a[5]  ^ ((~new_n471_ ^ ~\a[8] ) ^ ((new_n334_ & \a[8] ) | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] ))))))) ^ ((\a[5]  & ((new_n334_ & \a[8] ) | (~new_n334_ & ~\a[8] ) | ((~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))) & ((new_n334_ ^ \a[8] ) | (new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))) | (~new_n473_ & (~\a[5]  | ((~new_n334_ | ~\a[8] ) & (new_n334_ | \a[8] ) & ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))) | ((~new_n334_ ^ \a[8] ) & (~new_n335_ | ~\a[8] ) & (new_n337_ | (new_n335_ & \a[8] ) | (~new_n335_ & ~\a[8] )))) & (\a[5]  | ((new_n334_ ^ \a[8] ) ^ ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] )))))));
  assign new_n602_ = ((new_n473_ ^ ~new_n603_) | new_n582_ | ~\a[2] ) & ((new_n473_ & ~new_n603_) | (~new_n473_ & new_n603_) | (~new_n582_ & \a[2] )) & (~new_n604_ | new_n606_) & new_n607_ & (new_n604_ | ~new_n606_);
  assign new_n603_ = \a[5]  ^ ((new_n334_ ^ \a[8] ) ^ ((new_n335_ & \a[8] ) | (~new_n337_ & (~new_n335_ | ~\a[8] ) & (new_n335_ | \a[8] ))));
  assign new_n604_ = (~\a[2]  | (new_n480_ & ~new_n605_) | (~new_n480_ & new_n605_)) & ((\a[2]  & (~new_n480_ | new_n605_) & (new_n480_ | ~new_n605_)) | (~\a[2]  & (~new_n480_ ^ ~new_n605_)) | ((~new_n541_ | ~\a[2] ) & ((new_n541_ & \a[2] ) | (~new_n541_ & ~\a[2] ) | ((~new_n543_ | ~\a[2] ) & (new_n544_ | (~new_n543_ & ~\a[2] ) | (new_n543_ & \a[2] ))))));
  assign new_n605_ = \a[5]  ^ (new_n341_ ^ ~new_n479_);
  assign new_n606_ = \a[2]  ^ ((new_n477_ ^ \a[5] ) ^ ((new_n478_ & \a[5] ) | (~new_n480_ & (~new_n478_ | ~\a[5] ) & (new_n478_ | \a[5] ))));
  assign new_n607_ = ((new_n541_ & \a[2] ) | ((~new_n541_ | ~\a[2] ) & (new_n541_ | \a[2] ) & ((new_n543_ & \a[2] ) | ((~new_n543_ | ~\a[2] ) & (new_n543_ | \a[2] ) & ((new_n608_ & \a[2] ) | (~new_n609_ & (~new_n608_ | ~\a[2] ) & (new_n608_ | \a[2] )))))) | (\a[2]  ^ (new_n480_ ^ ~new_n605_))) & (((~new_n541_ | ~\a[2] ) & ((new_n541_ & \a[2] ) | (~new_n541_ & ~\a[2] ) | ((~new_n543_ | ~\a[2] ) & ((new_n543_ & \a[2] ) | (~new_n543_ & ~\a[2] ) | ((~new_n608_ | ~\a[2] ) & (new_n609_ | (new_n608_ & \a[2] ) | (~new_n608_ & ~\a[2] ))))))) | (\a[2]  & (~new_n480_ | new_n605_) & (new_n480_ | ~new_n605_)) | (~\a[2]  & (~new_n480_ ^ ~new_n605_))) & ((new_n541_ ^ \a[2] ) | (new_n543_ & \a[2] ) | ((~new_n543_ | ~\a[2] ) & (new_n543_ | \a[2] ) & ((new_n608_ & \a[2] ) | (~new_n609_ & (~new_n608_ | ~\a[2] ) & (new_n608_ | \a[2] ))))) & ((new_n541_ & \a[2] ) | (~new_n541_ & ~\a[2] ) | ((~new_n543_ | ~\a[2] ) & ((new_n543_ & \a[2] ) | (~new_n543_ & ~\a[2] ) | ((~new_n608_ | ~\a[2] ) & (new_n609_ | (new_n608_ & \a[2] ) | (~new_n608_ & ~\a[2] )))))) & ((~new_n543_ ^ \a[2] ) ^ ((new_n608_ & \a[2] ) | (~new_n609_ & (~new_n608_ | ~\a[2] ) & (new_n608_ | \a[2] )))) & new_n610_ & (new_n609_ ^ (new_n608_ ^ \a[2] ));
  assign new_n608_ = new_n484_ ^ ~new_n545_;
  assign new_n609_ = (~new_n546_ | new_n581_) & ((~new_n547_ & (new_n549_ | ~new_n580_)) | (new_n546_ & ~new_n581_) | (~new_n546_ & new_n581_));
  assign new_n610_ = (new_n612_ | new_n547_ | (new_n580_ & ((~new_n578_ & (new_n492_ | ~new_n516_) & (~new_n492_ | new_n516_)) | (~new_n611_ & (new_n578_ | (~new_n492_ & new_n516_) | (new_n492_ & ~new_n516_)) & (~new_n578_ | (~new_n492_ ^ new_n516_)))))) & (~new_n612_ | (~new_n547_ & (~new_n580_ | ((new_n578_ | (~new_n492_ & new_n516_) | (new_n492_ & ~new_n516_)) & (new_n611_ | (~new_n578_ & (new_n492_ | ~new_n516_) & (~new_n492_ | new_n516_)) | (new_n578_ & (new_n492_ ^ new_n516_))))))) & (~new_n580_ ^ ((~new_n578_ & (new_n492_ | ~new_n516_) & (~new_n492_ | new_n516_)) | (~new_n611_ & (new_n578_ | (~new_n492_ & new_n516_) | (new_n492_ & ~new_n516_)) & (~new_n578_ | (~new_n492_ ^ new_n516_))))) & new_n613_ & (new_n611_ ^ (~new_n578_ ^ (~new_n492_ ^ new_n516_)));
  assign new_n611_ = (~new_n550_ | new_n579_) & ((~new_n552_ & (new_n554_ | ~new_n577_)) | (new_n550_ & ~new_n579_) | (~new_n550_ & new_n579_));
  assign new_n612_ = ~new_n581_ ^ ((new_n487_ | (new_n517_ & (new_n489_ | (~new_n492_ & new_n516_)))) ^ (new_n485_ ^ ~new_n518_));
  assign new_n613_ = ((~new_n550_ ^ ~new_n579_) ^ (new_n552_ | (~new_n554_ & new_n577_))) & (~new_n554_ | new_n577_) & (new_n554_ | ~new_n577_) & (~new_n614_ | new_n615_) & new_n616_ & (new_n614_ | ~new_n615_);
  assign new_n614_ = (~new_n557_ | new_n576_) & ((~new_n558_ & (new_n560_ | ~new_n575_)) | (new_n557_ & ~new_n576_) | (~new_n557_ & new_n576_));
  assign new_n615_ = ~new_n556_ ^ (new_n498_ ^ ~new_n555_);
  assign new_n616_ = (~new_n619_ ^ (new_n558_ | (~new_n560_ & new_n575_))) & (~new_n560_ ^ ~new_n575_) & (~new_n617_ | new_n618_) & (new_n617_ | ~new_n618_) & ~new_n620_ & new_n621_;
  assign new_n617_ = (new_n563_ | ~new_n564_) & ((new_n563_ & ~new_n564_) | (~new_n563_ & new_n564_) | ((new_n565_ | ~new_n568_) & (new_n569_ | (~new_n565_ & new_n568_) | (new_n565_ & ~new_n568_))));
  assign new_n618_ = ~new_n562_ ^ (new_n506_ ^ ~new_n561_);
  assign new_n619_ = ~new_n576_ ^ ((new_n499_ ^ ~new_n500_) ^ ((new_n501_ & ~new_n502_) | ((new_n501_ | ~new_n502_) & (~new_n501_ | new_n502_) & ((~new_n503_ & new_n512_) | (~new_n506_ & (new_n503_ | ~new_n512_) & (~new_n503_ | new_n512_))))));
  assign new_n620_ = (new_n563_ ^ ~new_n564_) ^ ((~new_n565_ & new_n568_) | (~new_n569_ & (new_n565_ | ~new_n568_) & (~new_n565_ | new_n568_)));
  assign new_n621_ = (~new_n569_ | new_n622_) & (new_n569_ | ~new_n622_) & ~new_n623_ & ~new_n624_ & (new_n634_ | ~new_n635_) & (~new_n634_ | new_n635_) & new_n625_ & ~new_n636_;
  assign new_n622_ = (~new_n510_ ^ new_n511_) ^ (~\a[2]  ^ (new_n567_ & (~new_n60_ | ~new_n566_)));
  assign new_n623_ = (new_n571_ ^ (~\a[2]  ^ (new_n570_ & (~new_n63_ | ~new_n566_)))) ^ ((~new_n572_ & new_n573_) | (~new_n574_ & (new_n572_ | ~new_n573_) & (~new_n572_ | new_n573_)));
  assign new_n624_ = ~new_n574_ ^ (new_n572_ ^ ~new_n573_);
  assign new_n625_ = ~new_n627_ & (~new_n630_ | ~new_n631_ | ~new_n628_ | ~new_n629_) & new_n626_ & (~new_n632_ | ~new_n633_);
  assign new_n626_ = \a[0]  & \b[0] ;
  assign new_n627_ = ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[1]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[0]  | \a[0]  | ~\a[1] ) & (~\b[2]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[1]  | \a[0]  | ~\a[1] ) & (~\b[0]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )));
  assign new_n628_ = ~\a[27]  & ~\a[23]  & ~\a[24] ;
  assign new_n629_ = ~\a[21]  & ~\a[22]  & ~\a[25]  & ~\a[26]  & ~\a[17]  & ~\a[18]  & ~\a[19]  & ~\a[20] ;
  assign new_n630_ = ~\a[5]  & ~\a[6]  & ~\a[7]  & ~\a[8]  & ~\a[1]  & ~\a[2]  & ~\a[3]  & ~\a[4] ;
  assign new_n631_ = ~\a[11]  & ~\a[12]  & ~\a[15]  & ~\a[16]  & ~\a[9]  & ~\a[10]  & ~\a[13]  & ~\a[14] ;
  assign new_n632_ = ~\b[13]  & ~\b[14]  & ~\b[9]  & ~\b[10]  & ~\b[11]  & ~\b[12] ;
  assign new_n633_ = ~\b[5]  & ~\b[6]  & ~\b[7]  & ~\b[8]  & ~\b[2]  & ~\b[3]  & ~\b[1]  & ~\b[4] ;
  assign new_n634_ = \b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] );
  assign new_n635_ = \a[2]  ^ ((~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] ) & (~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )));
  assign new_n636_ = \a[2]  ? (((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[1]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[0]  & ~\a[0]  & \a[1] )) : ((\b[2]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[1]  & ~\a[0]  & \a[1] ) | (\b[0]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] ) & (~\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n637_ = ~new_n639_ ^ (~new_n638_ ^ (\a[5]  ^ ((\a[8]  & (~new_n428_ | new_n440_) & (new_n428_ | ~new_n440_)) | (((new_n522_ & \a[8] ) | (~new_n49_ & (~new_n522_ | ~\a[8] ) & (new_n522_ | \a[8] ))) & (~\a[8]  | (new_n428_ & ~new_n440_) | (~new_n428_ & new_n440_)) & (\a[8]  | (new_n428_ ^ ~new_n440_))))));
  assign new_n638_ = \a[17]  ^ ((\a[11]  & (new_n441_ | ~new_n442_) & (~new_n441_ | new_n442_)) | (~new_n428_ & (~\a[11]  | (~new_n441_ & new_n442_) | (new_n441_ & ~new_n442_)) & (\a[11]  | (~new_n441_ ^ new_n442_))));
  assign new_n639_ = new_n642_ ^ ((new_n641_ | (~new_n640_ & new_n448_)) ^ ((\a[20]  & (new_n640_ | ~new_n448_) & (~new_n640_ | new_n448_)) | (((new_n446_ & \a[20] ) | (~new_n432_ & (new_n446_ | \a[20] ) & (~new_n446_ | ~\a[20] ))) & (~\a[20]  | (~new_n640_ & new_n448_) | (new_n640_ & ~new_n448_)) & (\a[20]  | (~new_n640_ ^ new_n448_)))));
  assign new_n640_ = (~\a[23]  | (~new_n435_ & new_n438_) | (new_n435_ & ~new_n438_)) & (((~new_n434_ | ~\a[23] ) & (new_n415_ | (new_n434_ & \a[23] ) | (~new_n434_ & ~\a[23] ))) | (\a[23]  & (new_n435_ | ~new_n438_) & (~new_n435_ | new_n438_)) | (~\a[23]  & (new_n435_ ^ new_n438_)));
  assign new_n641_ = \a[23]  & (~new_n450_ | (~new_n449_ & (new_n435_ | ~new_n438_))) & (new_n450_ | new_n449_ | (~new_n435_ & new_n438_));
  assign new_n642_ = \a[14]  ^ ((\a[26]  & ((\a[27]  & \b[13] ) | (\b[14]  & (\a[26]  ^ \a[27] )))) | ((new_n449_ | (~new_n435_ & new_n438_)) & (~\a[26]  | ((~\a[27]  | ~\b[13] ) & (~\b[14]  | (~\a[26]  ^ \a[27] )))) & (\a[26]  | (\a[27]  & \b[14] ))));
endmodule


