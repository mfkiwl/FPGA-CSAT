// Benchmark "b17_C_sat" written by ABC on Fri Nov  4 11:02:37 2022

module b17_C_sat ( 
    P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
    DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
    DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
    DATAI_15_, DATAI_13_, DATAI_11_, DATAI_9_, DATAI_8_, DATAI_7_,
    DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_,
    HOLD, NA, BS16, READY1, READY2, P1_ADS_N_REG_SCAN_IN,
    P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
    P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
    P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
    P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
    P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
    P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
    P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN,
    P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN,
    P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN,
    P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN,
    P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN,
    P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN,
    P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN,
    P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN,
    P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN,
    P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
    P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN,
    P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_EBX_REG_31__SCAN_IN,
    P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
    P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN,
    P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
    P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN,
    P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
    P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN,
    P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN,
    P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN,
    P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN,
    P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN,
    P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
    P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN,
    P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
    P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN,
    P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
    P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN,
    P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
    P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
    P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
    P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
    P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
    P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
    P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
    P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
    P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN,
    P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN,
    P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_6__SCAN_IN,
    P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
    P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_3__SCAN_IN,
    P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
    P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
    P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_13__SCAN_IN,
    P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN,
    P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN,
    P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN,
    P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN,
    P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN,
    P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN,
    P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN,
    P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN,
    P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN,
    P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN,
    P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN,
    P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN,
    P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN,
    P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN,
    P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN,
    P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN,
    P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN,
    P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN,
    P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN,
    P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN,
    P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN,
    P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN,
    P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN,
    P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN,
    P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN,
    P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN,
    P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN,
    P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN,
    P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN,
    P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN,
    P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN,
    P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN,
    P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN,
    P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN,
    P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN,
    P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN,
    P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN,
    P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN,
    P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN,
    P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN,
    P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN,
    P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN,
    P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN,
    P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN,
    P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN,
    P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN,
    P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN,
    BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN,
    BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN,
    BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN,
    BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN,
    BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN,
    BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN,
    BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN,
    BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN,
    BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN,
    BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN,
    BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN,
    BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN,
    BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN,
    BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN,
    BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN,
    BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN,
    BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN,
    BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN,
    BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN,
    BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN,
    BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN,
    READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN,
    READY11_REG_SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
    P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
    P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN,
    P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN,
    P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN,
    P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
    P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
    P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
    P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN,
    P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN,
    P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN,
    P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN,
    P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN,
    P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN,
    P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN,
    P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN,
    P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN,
    P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN,
    P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN,
    P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN,
    P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN,
    P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN,
    P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN,
    P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN,
    P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN,
    P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN,
    P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN,
    P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN,
    P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN,
    P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN,
    P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN,
    P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN,
    P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN,
    P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN,
    P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN,
    P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN,
    P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN,
    P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN,
    P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN,
    P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN,
    P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN,
    P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN,
    P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN,
    P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN,
    P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN,
    P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN,
    P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN,
    P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN,
    P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN,
    P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN,
    P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN,
    P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN,
    P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN,
    P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN,
    P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN,
    P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN,
    P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN,
    P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN,
    P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN,
    P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN,
    P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN,
    P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN,
    P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN,
    P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN,
    P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN,
    P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN,
    P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN,
    P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN,
    P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN,
    P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN,
    P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN,
    P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN,
    P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN,
    P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN,
    P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN,
    P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN,
    P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN,
    P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN,
    P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN,
    P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN,
    P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN,
    P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN,
    P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN,
    P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN,
    P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN,
    P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN,
    P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN,
    P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN,
    P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN,
    P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN,
    P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN,
    P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
    P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
    P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
    P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
    P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
    P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
    P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN,
    P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN,
    P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN,
    P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN,
    P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN,
    P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN,
    P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN,
    P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN,
    P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN,
    P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN,
    P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
    P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
    P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
    P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
    P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
    P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
    P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
    P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
    P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
    P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
    P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
    P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
    P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
    P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
    P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
    P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
    P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_14__SCAN_IN,
    P3_LWORD_REG_13__SCAN_IN, P3_LWORD_REG_10__SCAN_IN,
    P3_LWORD_REG_9__SCAN_IN, P3_LWORD_REG_8__SCAN_IN,
    P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
    P3_LWORD_REG_1__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
    P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
    P3_UWORD_REG_10__SCAN_IN, P3_UWORD_REG_9__SCAN_IN,
    P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
    P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
    P3_UWORD_REG_1__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
    P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
    P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
    P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
    P3_DATAO_REG_31__SCAN_IN, P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN,
    P3_EAX_REG_2__SCAN_IN, P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN,
    P3_EAX_REG_5__SCAN_IN, P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN,
    P3_EAX_REG_8__SCAN_IN, P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN,
    P3_EAX_REG_11__SCAN_IN, P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
    P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN,
    P3_EAX_REG_17__SCAN_IN, P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
    P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN,
    P3_EAX_REG_23__SCAN_IN, P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
    P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN,
    P3_EAX_REG_29__SCAN_IN, P3_EAX_REG_30__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
    P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
    P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
    P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
    P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN,
    P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
    P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN,
    P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
    P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN,
    P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
    P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN,
    P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
    P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN,
    P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
    P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
    P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
    P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
    P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
    P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
    P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
    P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
    P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
    P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
    P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
    P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
    P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
    P3_BYTEENABLE_REG_3__SCAN_IN, P3_FLUSH_REG_SCAN_IN,
    P3_MORE_REG_SCAN_IN, P3_STATEBS16_REG_SCAN_IN,
    P3_REQUESTPENDING_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN,
    P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
    P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN,
    P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN,
    P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN,
    P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN,
    P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN,
    P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN,
    P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN,
    P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN,
    P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN,
    P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN,
    P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN,
    P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN,
    P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN,
    P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN,
    P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN,
    P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN,
    P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN,
    P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN,
    P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN,
    P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN,
    P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN,
    P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN,
    P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN,
    P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN,
    P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN,
    P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN,
    P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN,
    P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN,
    P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN,
    P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN,
    P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN,
    P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN,
    P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN,
    P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN,
    P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN,
    P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN,
    P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN,
    P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN,
    P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN,
    P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN,
    P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN,
    P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN,
    P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN,
    P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN,
    P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN,
    P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN,
    P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN,
    P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN,
    P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN,
    P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN,
    P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN,
    P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN,
    P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN,
    P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN,
    P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN,
    P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN,
    P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN,
    P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN,
    P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN,
    P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN,
    P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN,
    P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN,
    P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN,
    P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN,
    P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN,
    P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN,
    P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN,
    P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN,
    P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN,
    P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN,
    P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN,
    P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN,
    P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN,
    P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN,
    P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN,
    P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN,
    P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN,
    P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN,
    P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN,
    P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN,
    P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN,
    P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN,
    P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN,
    P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN,
    P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN,
    P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN,
    P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN,
    P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN,
    P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN,
    P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN,
    P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN,
    P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN,
    P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN,
    P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN,
    P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN,
    P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN,
    P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN,
    P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN,
    P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN,
    P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
    P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
    P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
    P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
    P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
    P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
    P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN,
    P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN,
    P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN,
    P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN,
    P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN,
    P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN,
    P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN,
    P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN,
    P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN,
    P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN,
    P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
    P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
    P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
    P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
    P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
    P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
    P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
    P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
    P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
    P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
    P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
    P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
    P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
    P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
    P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
    P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
    P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
    P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_10__SCAN_IN,
    P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
    P2_LWORD_REG_3__SCAN_IN, P2_LWORD_REG_2__SCAN_IN,
    P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_7__SCAN_IN,
    P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
    P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_1__SCAN_IN,
    P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
    P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
    P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
    P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
    P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
    P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
    P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
    P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
    P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN,
    P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
    P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN,
    P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
    P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN,
    P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
    P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
    P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
    P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
    P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
    P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN,
    P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
    P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN,
    P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
    P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN,
    P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
    P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN,
    P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
    P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN,
    P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
    P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
    P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
    P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
    P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
    P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
    P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
    P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
    P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
    P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
    P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
    P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
    P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
    P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
    P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
    P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
    P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
    P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
    P1_BE_N_REG_3__SCAN_IN, P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
    P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
    P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
    P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
    P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
    P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
    P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
    P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
    P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
    P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
    P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
    P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
    P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
    P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
    P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
    P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
    P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
    P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
    P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
    P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN,
    P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN,
    P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN,
    P1_DATAWIDTH_REG_30__SCAN_IN, P1_STATE2_REG_3__SCAN_IN,
    P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN,
    P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN,
    P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN,
    P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN,
    P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN,
    P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN,
    P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN,
    P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN,
    P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN,
    P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN,
    P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN,
    P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN,
    P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN,
    P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN,
    P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN,
    P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN,
    P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN,
    P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN,
    P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN,
    P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN,
    P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN,
    P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN,
    P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN,
    P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN,
    P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN,
    P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN,
    P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN,
    P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN,
    P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN,
    P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN,
    P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN,
    P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN,
    P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN,
    P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN,
    P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN,
    P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN,
    P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN,
    P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN,
    P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN,
    P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN,
    P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN,
    P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN,
    P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN,
    P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN,
    P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN,
    P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN,
    P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN,
    P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN,
    sat  );
  input  P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_,
    DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
    DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
    DATAI_16_, DATAI_15_, DATAI_13_, DATAI_11_, DATAI_9_, DATAI_8_,
    DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
    DATAI_0_, HOLD, NA, BS16, READY1, READY2, P1_ADS_N_REG_SCAN_IN,
    P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
    P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
    P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
    P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
    P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
    P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
    P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN,
    P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN,
    P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN,
    P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN,
    P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN,
    P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN,
    P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN,
    P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN,
    P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN,
    P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
    P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN,
    P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_EBX_REG_31__SCAN_IN,
    P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
    P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN,
    P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
    P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN,
    P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
    P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN,
    P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN,
    P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN,
    P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN,
    P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN,
    P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
    P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN,
    P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
    P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN,
    P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
    P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN,
    P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
    P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
    P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
    P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
    P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
    P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
    P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
    P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
    P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN,
    P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN,
    P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_6__SCAN_IN,
    P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
    P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_3__SCAN_IN,
    P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
    P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
    P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_13__SCAN_IN,
    P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN,
    P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN,
    P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN,
    P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN,
    P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN,
    P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN,
    P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN,
    P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN,
    P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN,
    P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN,
    P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN,
    P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN,
    P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN,
    P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN,
    P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN,
    P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN,
    P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN,
    P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN,
    P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN,
    P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN,
    P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN,
    P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN,
    P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN,
    P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN,
    P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN,
    P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN,
    P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN,
    P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN,
    P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN,
    P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN,
    P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN,
    P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN,
    P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN,
    P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN,
    P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN,
    P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN,
    P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN,
    P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN,
    P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN,
    P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN,
    P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN,
    P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN,
    P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN,
    P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN,
    P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN,
    P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN,
    P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN,
    BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN,
    BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN,
    BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN,
    BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN,
    BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN,
    BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN,
    BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN,
    BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN,
    BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN,
    BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN,
    BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN,
    BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN,
    BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN,
    BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN,
    BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN,
    BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN,
    BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN,
    BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN,
    BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN,
    BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN,
    BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN,
    READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN,
    READY11_REG_SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
    P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
    P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN,
    P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN,
    P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN,
    P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
    P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
    P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
    P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN,
    P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN,
    P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN,
    P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN,
    P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN,
    P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN,
    P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN,
    P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN,
    P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN,
    P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN,
    P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN,
    P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN,
    P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN,
    P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN,
    P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN,
    P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN,
    P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN,
    P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN,
    P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN,
    P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN,
    P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN,
    P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN,
    P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN,
    P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN,
    P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN,
    P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN,
    P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN,
    P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN,
    P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN,
    P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN,
    P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN,
    P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN,
    P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN,
    P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN,
    P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN,
    P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN,
    P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN,
    P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN,
    P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN,
    P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN,
    P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN,
    P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN,
    P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN,
    P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN,
    P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN,
    P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN,
    P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN,
    P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN,
    P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN,
    P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN,
    P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN,
    P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN,
    P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN,
    P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN,
    P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN,
    P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN,
    P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN,
    P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN,
    P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN,
    P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN,
    P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN,
    P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN,
    P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN,
    P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN,
    P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN,
    P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN,
    P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN,
    P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN,
    P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN,
    P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN,
    P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN,
    P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN,
    P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN,
    P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN,
    P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN,
    P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN,
    P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN,
    P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN,
    P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN,
    P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN,
    P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN,
    P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN,
    P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN,
    P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
    P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
    P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
    P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
    P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
    P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
    P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN,
    P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN,
    P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN,
    P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN,
    P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN,
    P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN,
    P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN,
    P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN,
    P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN,
    P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN,
    P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
    P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
    P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
    P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
    P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
    P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
    P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
    P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
    P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
    P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
    P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
    P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
    P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
    P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
    P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
    P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
    P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_14__SCAN_IN,
    P3_LWORD_REG_13__SCAN_IN, P3_LWORD_REG_10__SCAN_IN,
    P3_LWORD_REG_9__SCAN_IN, P3_LWORD_REG_8__SCAN_IN,
    P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
    P3_LWORD_REG_1__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
    P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
    P3_UWORD_REG_10__SCAN_IN, P3_UWORD_REG_9__SCAN_IN,
    P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
    P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
    P3_UWORD_REG_1__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
    P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
    P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
    P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
    P3_DATAO_REG_31__SCAN_IN, P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN,
    P3_EAX_REG_2__SCAN_IN, P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN,
    P3_EAX_REG_5__SCAN_IN, P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN,
    P3_EAX_REG_8__SCAN_IN, P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN,
    P3_EAX_REG_11__SCAN_IN, P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
    P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN,
    P3_EAX_REG_17__SCAN_IN, P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
    P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN,
    P3_EAX_REG_23__SCAN_IN, P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
    P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN,
    P3_EAX_REG_29__SCAN_IN, P3_EAX_REG_30__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
    P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
    P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
    P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
    P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN,
    P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
    P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN,
    P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
    P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN,
    P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
    P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN,
    P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
    P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN,
    P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
    P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
    P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
    P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
    P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
    P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
    P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
    P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
    P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
    P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
    P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
    P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
    P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
    P3_BYTEENABLE_REG_3__SCAN_IN, P3_FLUSH_REG_SCAN_IN,
    P3_MORE_REG_SCAN_IN, P3_STATEBS16_REG_SCAN_IN,
    P3_REQUESTPENDING_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN,
    P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
    P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN,
    P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN,
    P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN,
    P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN,
    P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN,
    P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN,
    P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN,
    P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN,
    P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN,
    P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN,
    P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN,
    P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN,
    P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN,
    P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN,
    P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN,
    P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN,
    P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN,
    P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN,
    P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN,
    P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN,
    P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN,
    P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN,
    P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN,
    P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN,
    P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN,
    P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN,
    P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN,
    P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN,
    P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN,
    P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN,
    P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN,
    P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN,
    P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN,
    P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN,
    P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN,
    P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN,
    P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN,
    P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN,
    P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN,
    P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN,
    P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN,
    P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN,
    P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN,
    P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN,
    P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN,
    P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN,
    P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN,
    P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN,
    P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN,
    P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN,
    P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN,
    P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN,
    P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN,
    P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN,
    P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN,
    P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN,
    P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN,
    P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN,
    P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN,
    P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN,
    P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN,
    P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN,
    P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN,
    P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN,
    P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN,
    P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN,
    P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN,
    P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN,
    P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN,
    P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN,
    P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN,
    P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN,
    P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN,
    P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN,
    P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN,
    P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN,
    P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN,
    P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN,
    P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN,
    P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN,
    P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN,
    P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN,
    P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN,
    P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN,
    P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN,
    P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN,
    P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN,
    P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN,
    P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN,
    P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN,
    P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN,
    P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN,
    P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN,
    P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN,
    P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN,
    P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN,
    P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN,
    P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN,
    P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN,
    P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
    P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
    P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
    P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
    P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
    P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
    P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN,
    P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN,
    P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN,
    P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN,
    P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN,
    P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN,
    P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN,
    P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN,
    P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN,
    P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN,
    P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
    P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
    P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
    P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
    P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
    P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
    P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
    P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
    P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
    P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
    P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
    P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
    P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
    P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
    P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
    P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
    P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
    P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_10__SCAN_IN,
    P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
    P2_LWORD_REG_3__SCAN_IN, P2_LWORD_REG_2__SCAN_IN,
    P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_7__SCAN_IN,
    P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
    P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_1__SCAN_IN,
    P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
    P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
    P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
    P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
    P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
    P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
    P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
    P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
    P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN,
    P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
    P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN,
    P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
    P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN,
    P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
    P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
    P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
    P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
    P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
    P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN,
    P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
    P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN,
    P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
    P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN,
    P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
    P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN,
    P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
    P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN,
    P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
    P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
    P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
    P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
    P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
    P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
    P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
    P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
    P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
    P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
    P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
    P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
    P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
    P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
    P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
    P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
    P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
    P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
    P1_BE_N_REG_3__SCAN_IN, P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
    P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
    P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
    P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
    P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
    P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
    P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
    P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
    P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
    P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
    P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
    P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
    P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
    P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
    P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
    P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
    P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
    P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
    P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
    P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN,
    P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN,
    P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN,
    P1_DATAWIDTH_REG_30__SCAN_IN, P1_STATE2_REG_3__SCAN_IN,
    P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN,
    P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN,
    P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN,
    P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN,
    P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN,
    P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN,
    P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN,
    P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN,
    P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN,
    P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN,
    P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN,
    P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN,
    P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN,
    P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN,
    P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN,
    P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN,
    P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN,
    P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN,
    P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN,
    P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN,
    P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN,
    P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN,
    P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN,
    P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN,
    P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN,
    P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN,
    P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN,
    P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN,
    P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN,
    P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN,
    P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN,
    P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN,
    P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN,
    P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN,
    P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN,
    P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN,
    P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN,
    P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN,
    P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN,
    P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN,
    P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN,
    P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN,
    P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN,
    P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN,
    P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN,
    P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN,
    P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN,
    P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output sat;
  wire new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_,
    new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_,
    new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_,
    new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_,
    new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_,
    new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_,
    new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_,
    new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_,
    new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_,
    new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_,
    new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_,
    new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_,
    new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_,
    new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_,
    new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_,
    new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_,
    new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_,
    new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_,
    new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_,
    new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_,
    new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_,
    new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_,
    new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_,
    new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_,
    new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_,
    new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_,
    new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_,
    new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_,
    new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_,
    new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_,
    new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_,
    new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_,
    new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_,
    new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_,
    new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_,
    new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_,
    new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_,
    new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_,
    new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_,
    new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_,
    new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_,
    new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_,
    new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_,
    new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_,
    new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_,
    new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_,
    new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_,
    new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_,
    new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_,
    new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_,
    new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_,
    new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_,
    new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_,
    new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_,
    new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_,
    new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_,
    new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_,
    new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_,
    new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_,
    new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_,
    new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_,
    new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_,
    new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_,
    new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_,
    new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_,
    new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_,
    new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_,
    new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_,
    new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_,
    new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_,
    new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_,
    new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_,
    new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_,
    new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_,
    new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_,
    new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_,
    new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_,
    new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_,
    new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_,
    new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_,
    new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_,
    new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_,
    new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_,
    new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_,
    new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_,
    new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_,
    new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_,
    new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_,
    new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_,
    new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_,
    new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_,
    new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_,
    new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_,
    new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_,
    new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_,
    new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_,
    new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_,
    new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_,
    new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_,
    new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_, new_n3276_,
    new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_,
    new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_,
    new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_,
    new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_,
    new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_,
    new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_,
    new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_,
    new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_,
    new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_,
    new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_,
    new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_,
    new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_,
    new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_,
    new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_,
    new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_,
    new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_,
    new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_,
    new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_,
    new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_,
    new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_,
    new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_,
    new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_,
    new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_,
    new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_,
    new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_,
    new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_,
    new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_,
    new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_,
    new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_,
    new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_,
    new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_,
    new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_,
    new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_,
    new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_,
    new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_,
    new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_,
    new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_,
    new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_,
    new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_,
    new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_,
    new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_,
    new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_,
    new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_,
    new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_,
    new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_,
    new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_,
    new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_,
    new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_,
    new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_,
    new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_,
    new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_,
    new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_,
    new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_,
    new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_,
    new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_,
    new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_,
    new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_,
    new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_,
    new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_,
    new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_,
    new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_,
    new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_,
    new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_,
    new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_,
    new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_,
    new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_,
    new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_, new_n3678_,
    new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_,
    new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_,
    new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_,
    new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_,
    new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_,
    new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_,
    new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_,
    new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_, new_n3726_,
    new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_, new_n3732_,
    new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_, new_n3738_,
    new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_,
    new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_,
    new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_,
    new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_,
    new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_,
    new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_, new_n3774_,
    new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_,
    new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_,
    new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_,
    new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_,
    new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_,
    new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_,
    new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_,
    new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_,
    new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_,
    new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_,
    new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_,
    new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_,
    new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_,
    new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_,
    new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_,
    new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_,
    new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_,
    new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_,
    new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_,
    new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_,
    new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_,
    new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_,
    new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_,
    new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_,
    new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_,
    new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_,
    new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_,
    new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_,
    new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_,
    new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_,
    new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_,
    new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_,
    new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_, new_n3972_,
    new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_, new_n3978_,
    new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_, new_n3984_,
    new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_, new_n3990_,
    new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_, new_n3996_,
    new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_, new_n4002_,
    new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_, new_n4008_,
    new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_, new_n4014_,
    new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_,
    new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_,
    new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_,
    new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_,
    new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_,
    new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_,
    new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_,
    new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_,
    new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_,
    new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_,
    new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_,
    new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_,
    new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_,
    new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_,
    new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_,
    new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_,
    new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_,
    new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_,
    new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_, new_n4128_,
    new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_, new_n4134_,
    new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_, new_n4140_,
    new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_,
    new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_,
    new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_,
    new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_,
    new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_,
    new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_,
    new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_,
    new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_,
    new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_,
    new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_,
    new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_,
    new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_,
    new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_,
    new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_,
    new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_,
    new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_,
    new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_,
    new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_,
    new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_,
    new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_,
    new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_,
    new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_,
    new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_,
    new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_,
    new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_,
    new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_,
    new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_,
    new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_,
    new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_,
    new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_,
    new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_,
    new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_,
    new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_,
    new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_,
    new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_,
    new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_,
    new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_,
    new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_,
    new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_,
    new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_,
    new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_,
    new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_,
    new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_,
    new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_,
    new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_,
    new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_,
    new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_,
    new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_,
    new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_,
    new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_,
    new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_,
    new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_,
    new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_,
    new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_,
    new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_,
    new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_,
    new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_,
    new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_,
    new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_,
    new_n4513_, new_n4514_;
  assign sat = ~new_n1304_ & new_n1793_ & (~new_n4509_ | ((new_n4508_ | (new_n4514_ ^ P2_INSTADDRPOINTER_REG_30__SCAN_IN)) & new_n4420_ & (~new_n4508_ | (new_n4514_ & P2_INSTADDRPOINTER_REG_30__SCAN_IN) | (~new_n4514_ & ~P2_INSTADDRPOINTER_REG_30__SCAN_IN))));
  assign new_n1304_ = (new_n1750_ | ((~new_n1729_ | (~new_n1305_ & new_n1749_)) & (new_n1730_ | new_n1743_))) & new_n1758_ & (~new_n1750_ | (new_n1729_ & (new_n1305_ | ~new_n1749_)) | (~new_n1730_ & ~new_n1743_));
  assign new_n1305_ = new_n1711_ & (new_n1728_ | (~new_n1306_ & (~new_n1526_ | (~new_n1308_ & ~new_n1630_) | (new_n1308_ & new_n1630_))));
  assign new_n1306_ = ~new_n1307_ & ((new_n1701_ & new_n1702_) | ((new_n1701_ | new_n1702_) & ((new_n1705_ & ~new_n1706_) | ((new_n1705_ | ~new_n1706_) & (new_n1708_ | (~new_n1637_ & ~new_n1710_))))));
  assign new_n1307_ = ~new_n1526_ & (~new_n1308_ ^ new_n1630_);
  assign new_n1308_ = (~new_n1509_ | ((~new_n1510_ | ~new_n1309_ | new_n1520_) & (~new_n1497_ | ~new_n1316_ | ~new_n1322_)) | ((new_n1515_ | ~new_n1316_ | ~new_n1322_) & ((~new_n1497_ & new_n1515_) | ~new_n1316_ | new_n1322_ | (new_n1497_ & ~new_n1515_)))) & (new_n1515_ | ~new_n1316_ | ~new_n1322_ | new_n1322_ | (new_n1497_ & ~new_n1515_));
  assign new_n1309_ = new_n1486_ & ~new_n1491_ & new_n1310_ & new_n1481_;
  assign new_n1310_ = ~new_n1476_ & new_n1466_ & new_n1459_ & new_n1311_ & ~new_n1471_;
  assign new_n1311_ = new_n1422_ & ~new_n1454_ & new_n1428_ & ~new_n1448_ & new_n1436_ & ~new_n1443_ & new_n1312_ & new_n1442_;
  assign new_n1312_ = P2_INSTQUEUE_REG_0__6__SCAN_IN & new_n1419_ & ~new_n1420_ & (new_n1313_ | (~new_n1408_ & (~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_))));
  assign new_n1313_ = new_n1314_ & (~new_n1405_ | (new_n1407_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_))));
  assign new_n1314_ = new_n1315_ & P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign new_n1315_ = new_n1316_ & ~new_n1322_;
  assign new_n1316_ = new_n1317_ & P2_STATE2_REG_0__SCAN_IN;
  assign new_n1317_ = new_n1320_ & new_n1321_ & new_n1318_ & new_n1319_;
  assign new_n1318_ = (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_12__6__SCAN_IN : ~P2_INSTQUEUE_REG_4__6__SCAN_IN)) & (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_1__6__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_9__6__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1319_ = ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_11__6__SCAN_IN : ~P2_INSTQUEUE_REG_3__6__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & ((~P2_INSTQUEUE_REG_0__6__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_8__6__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1320_ = ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_14__6__SCAN_IN : ~P2_INSTQUEUE_REG_6__6__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_10__6__SCAN_IN : ~P2_INSTQUEUE_REG_2__6__SCAN_IN));
  assign new_n1321_ = ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_15__6__SCAN_IN : ~P2_INSTQUEUE_REG_7__6__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_13__6__SCAN_IN : ~P2_INSTQUEUE_REG_5__6__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1322_ = new_n1325_ & new_n1326_ & new_n1323_ & new_n1324_;
  assign new_n1323_ = ((~P2_INSTQUEUE_REG_0__1__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_8__1__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_11__1__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_3__1__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1324_ = (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_1__1__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_9__1__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN)) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_12__1__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_4__1__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1325_ = (~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_15__1__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_7__1__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN)) & ((~P2_INSTQUEUE_REG_5__1__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_13__1__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1326_ = ((~P2_INSTQUEUE_REG_2__1__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_10__1__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_14__1__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_6__1__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1327_ = ((new_n1382_ & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN & (~new_n1328_ | ~new_n1365_))) ^ (~new_n1379_ | (~new_n1373_ & P2_INSTADDRPOINTER_REG_3__SCAN_IN));
  assign new_n1328_ = ~new_n1329_ & ~new_n1355_ & ~new_n1357_;
  assign new_n1329_ = ~new_n1322_ & new_n1340_ & ~new_n1345_ & (((new_n1330_ ^ new_n1317_) & (new_n1330_ | new_n1350_)) | new_n1335_ | (~new_n1350_ & (new_n1330_ | ~new_n1317_)));
  assign new_n1330_ = new_n1333_ & new_n1334_ & new_n1331_ & new_n1332_;
  assign new_n1331_ = (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_1__5__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_9__5__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN)) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_12__5__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_4__5__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1332_ = ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_11__5__SCAN_IN : ~P2_INSTQUEUE_REG_3__5__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & ((~P2_INSTQUEUE_REG_0__5__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_8__5__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1333_ = ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_14__5__SCAN_IN : ~P2_INSTQUEUE_REG_6__5__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_10__5__SCAN_IN : ~P2_INSTQUEUE_REG_2__5__SCAN_IN));
  assign new_n1334_ = ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_15__5__SCAN_IN : ~P2_INSTQUEUE_REG_7__5__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_13__5__SCAN_IN : ~P2_INSTQUEUE_REG_5__5__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1335_ = new_n1338_ & new_n1339_ & new_n1336_ & new_n1337_;
  assign new_n1336_ = (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_12__7__SCAN_IN : ~P2_INSTQUEUE_REG_4__7__SCAN_IN)) & (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_1__7__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_9__7__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1337_ = ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_11__7__SCAN_IN : ~P2_INSTQUEUE_REG_3__7__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & ((~P2_INSTQUEUE_REG_0__7__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_8__7__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1338_ = ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_14__7__SCAN_IN : ~P2_INSTQUEUE_REG_6__7__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_10__7__SCAN_IN : ~P2_INSTQUEUE_REG_2__7__SCAN_IN));
  assign new_n1339_ = ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_15__7__SCAN_IN : ~P2_INSTQUEUE_REG_7__7__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_13__7__SCAN_IN : ~P2_INSTQUEUE_REG_5__7__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1340_ = P2_STATE2_REG_0__SCAN_IN & (~new_n1343_ | ~new_n1344_ | ~new_n1341_ | ~new_n1342_);
  assign new_n1341_ = ((~P2_INSTQUEUE_REG_0__0__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_8__0__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_11__0__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_3__0__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1342_ = (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_1__0__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_9__0__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN)) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_12__0__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_4__0__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1343_ = (~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_15__0__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_7__0__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN)) & ((~P2_INSTQUEUE_REG_5__0__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_13__0__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1344_ = ((~P2_INSTQUEUE_REG_2__0__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_10__0__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_14__0__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_6__0__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1345_ = new_n1348_ & new_n1349_ & new_n1346_ & new_n1347_;
  assign new_n1346_ = (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_12__3__SCAN_IN : ~P2_INSTQUEUE_REG_4__3__SCAN_IN)) & (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_1__3__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_9__3__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1347_ = ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_11__3__SCAN_IN : ~P2_INSTQUEUE_REG_3__3__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & ((~P2_INSTQUEUE_REG_0__3__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_8__3__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1348_ = (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_10__3__SCAN_IN : ~P2_INSTQUEUE_REG_2__3__SCAN_IN)) & (~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_14__3__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_6__3__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1349_ = ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_15__3__SCAN_IN : ~P2_INSTQUEUE_REG_7__3__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_13__3__SCAN_IN : ~P2_INSTQUEUE_REG_5__3__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1350_ = new_n1353_ & new_n1354_ & new_n1351_ & new_n1352_;
  assign new_n1351_ = (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_12__4__SCAN_IN : ~P2_INSTQUEUE_REG_4__4__SCAN_IN)) & (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_1__4__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_9__4__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1352_ = ((~P2_INSTQUEUE_REG_0__4__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_8__4__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_11__4__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_3__4__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1353_ = ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_14__4__SCAN_IN : ~P2_INSTQUEUE_REG_6__4__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_10__4__SCAN_IN : ~P2_INSTQUEUE_REG_2__4__SCAN_IN));
  assign new_n1354_ = ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_15__4__SCAN_IN : ~P2_INSTQUEUE_REG_7__4__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & ((~P2_INSTQUEUE_REG_5__4__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_13__4__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1355_ = ((~new_n1330_ & new_n1317_) | (new_n1330_ & ~new_n1317_) | ~new_n1350_ | ~new_n1356_) & new_n1322_ & new_n1340_;
  assign new_n1356_ = (~new_n1338_ | ~new_n1339_ | ~new_n1336_ | ~new_n1337_) & (~new_n1346_ | ~new_n1347_ | ~new_n1348_ | ~new_n1349_);
  assign new_n1357_ = P2_STATE2_REG_0__SCAN_IN & new_n1364_ & new_n1359_ & new_n1358_ & new_n1330_ & ~new_n1317_;
  assign new_n1358_ = new_n1338_ & new_n1339_ & new_n1336_ & new_n1337_ & new_n1351_ & new_n1352_ & new_n1353_ & new_n1354_;
  assign new_n1359_ = new_n1348_ & new_n1349_ & new_n1346_ & new_n1347_ & new_n1360_ & new_n1361_ & new_n1362_ & new_n1363_;
  assign new_n1360_ = (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_12__2__SCAN_IN : ~P2_INSTQUEUE_REG_4__2__SCAN_IN)) & (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_9__2__SCAN_IN : ~P2_INSTQUEUE_REG_1__2__SCAN_IN));
  assign new_n1361_ = ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_11__2__SCAN_IN : ~P2_INSTQUEUE_REG_3__2__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & ((~P2_INSTQUEUE_REG_0__2__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_8__2__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1362_ = ((~P2_INSTQUEUE_REG_2__2__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_10__2__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_14__2__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (~P2_INSTQUEUE_REG_6__2__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1363_ = ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_15__2__SCAN_IN : ~P2_INSTQUEUE_REG_7__2__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_13__2__SCAN_IN : ~P2_INSTQUEUE_REG_5__2__SCAN_IN) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1364_ = new_n1325_ & new_n1326_ & new_n1323_ & new_n1324_ & new_n1341_ & new_n1342_ & new_n1343_ & new_n1344_;
  assign new_n1365_ = ~new_n1372_ & ~new_n1366_ & ~new_n1369_ & ~new_n1371_;
  assign new_n1366_ = new_n1322_ & new_n1368_ & ((~new_n1367_ & (new_n1335_ | new_n1317_ | new_n1330_ | ~new_n1350_)) | (new_n1350_ ? (new_n1317_ & new_n1367_) : new_n1335_) | ((new_n1330_ | ~new_n1317_) & (~new_n1345_ | (~new_n1330_ & new_n1367_))));
  assign new_n1367_ = new_n1362_ & new_n1363_ & new_n1360_ & new_n1361_;
  assign new_n1368_ = P2_STATE2_REG_0__SCAN_IN & new_n1343_ & new_n1344_ & new_n1341_ & new_n1342_;
  assign new_n1369_ = ~new_n1322_ & P2_STATE2_REG_0__SCAN_IN & (new_n1370_ | (new_n1345_ & (~new_n1358_ | ~new_n1330_ | new_n1317_)));
  assign new_n1370_ = new_n1343_ & new_n1344_ & new_n1341_ & new_n1342_;
  assign new_n1371_ = new_n1340_ & (~new_n1367_ | (new_n1356_ & new_n1367_ & ~new_n1317_ & ~new_n1330_ & new_n1350_));
  assign new_n1372_ = ~new_n1330_ & new_n1317_ & new_n1322_ & new_n1368_;
  assign new_n1373_ = (new_n1374_ | ~P2_STATE2_REG_0__SCAN_IN) & ~new_n1376_ & (~new_n1375_ | ~P2_STATE2_REG_0__SCAN_IN);
  assign new_n1374_ = (new_n1335_ | new_n1317_ | new_n1330_ | ~new_n1350_ | ~new_n1370_ | ~new_n1345_ | new_n1367_) & (~new_n1345_ | ~new_n1367_ | ~new_n1330_ | new_n1335_ | ~new_n1322_ | new_n1317_ | ~new_n1370_);
  assign new_n1375_ = new_n1359_ & new_n1330_ & ~new_n1335_ & ~new_n1350_ & new_n1317_ & new_n1364_;
  assign new_n1376_ = new_n1322_ & new_n1340_ & ~new_n1378_ & new_n1330_ & new_n1377_ & new_n1350_ & new_n1356_;
  assign new_n1377_ = new_n1320_ & new_n1321_ & new_n1318_ & new_n1319_ & new_n1360_ & new_n1361_ & new_n1362_ & new_n1363_;
  assign new_n1378_ = P2_STATE_REG_2__SCAN_IN ^ ~P2_STATE_REG_1__SCAN_IN;
  assign new_n1379_ = (~new_n1380_ | ~P2_REIP_REG_3__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_3__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_3__SCAN_IN);
  assign new_n1380_ = new_n1330_ & new_n1377_ & new_n1350_ & new_n1356_ & ~new_n1322_ & new_n1340_;
  assign new_n1381_ = ~new_n1322_ & new_n1340_ & new_n1359_ & new_n1358_ & new_n1330_ & ~new_n1317_;
  assign new_n1382_ = ~P2_STATE2_REG_1__SCAN_IN & ~P2_STATE2_REG_0__SCAN_IN;
  assign new_n1383_ = (~new_n1384_ | (~new_n1373_ & P2_INSTADDRPOINTER_REG_2__SCAN_IN)) & (~new_n1385_ | (P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & (~new_n1328_ | ~new_n1365_)));
  assign new_n1384_ = (~new_n1380_ | ~P2_REIP_REG_2__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_2__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_2__SCAN_IN);
  assign new_n1385_ = ~P2_STATE2_REG_1__SCAN_IN & (P2_STATE2_REG_0__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  assign new_n1386_ = new_n1384_ & (new_n1373_ | ~P2_INSTADDRPOINTER_REG_2__SCAN_IN) & new_n1385_ & (~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | (new_n1328_ & new_n1365_));
  assign new_n1387_ = (new_n1398_ | new_n1390_ | (new_n1328_ & new_n1388_) | (~new_n1391_ & new_n1392_)) & ((~new_n1401_ & new_n1402_) | (new_n1398_ & (new_n1390_ | (new_n1328_ & new_n1388_) | (~new_n1391_ & new_n1392_))));
  assign new_n1388_ = ~new_n1366_ & ~new_n1369_ & ~new_n1371_ & ~new_n1372_ & new_n1389_ & (~new_n1375_ | ~P2_STATE2_REG_0__SCAN_IN);
  assign new_n1389_ = (~new_n1382_ | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (new_n1322_ | ~new_n1340_ | ~new_n1359_ | ~new_n1358_ | ~new_n1330_ | new_n1317_);
  assign new_n1390_ = ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & new_n1389_ & (~new_n1375_ | ~P2_STATE2_REG_0__SCAN_IN);
  assign new_n1391_ = P2_INSTADDRPOINTER_REG_0__SCAN_IN & ((~new_n1374_ & P2_STATE2_REG_0__SCAN_IN) | new_n1376_ | (new_n1375_ & P2_STATE2_REG_0__SCAN_IN));
  assign new_n1392_ = ~new_n1394_ & new_n1396_ & (~new_n1381_ | ~P2_EBX_REG_0__SCAN_IN) & (new_n1393_ | new_n1395_);
  assign new_n1393_ = (new_n1367_ | (~new_n1335_ & ~new_n1317_ & ~new_n1330_ & new_n1350_)) & (new_n1350_ ? (~new_n1317_ | ~new_n1367_) : ~new_n1335_) & ((~new_n1330_ & new_n1317_) | (new_n1345_ & (new_n1330_ | ~new_n1367_)));
  assign new_n1394_ = ((~new_n1345_ & (((new_n1330_ ^ new_n1317_) & (new_n1330_ | new_n1350_)) | new_n1335_ | (~new_n1350_ & (new_n1330_ | ~new_n1317_)))) | new_n1370_ | (new_n1345_ & (~new_n1330_ | new_n1317_ | ~new_n1335_ | ~new_n1350_))) & P2_STATE2_REG_0__SCAN_IN & ((new_n1330_ & ~new_n1317_ & new_n1335_ & new_n1350_) | ~new_n1322_ | (~new_n1330_ & new_n1317_));
  assign new_n1395_ = (~new_n1322_ | ~new_n1370_ | ~P2_STATE2_REG_0__SCAN_IN) & (~P2_REIP_REG_0__SCAN_IN | ~new_n1330_ | ~new_n1377_ | ~new_n1350_ | ~new_n1356_ | new_n1322_ | new_n1370_ | ~P2_STATE2_REG_0__SCAN_IN);
  assign new_n1396_ = (~new_n1340_ | (new_n1367_ & (~new_n1356_ | ~new_n1367_ | new_n1317_ | new_n1330_ | ~new_n1350_))) & new_n1397_ & (((new_n1330_ | ~new_n1317_) & (~new_n1330_ | new_n1317_) & new_n1350_ & new_n1356_) | ~new_n1322_ | ~new_n1340_);
  assign new_n1397_ = P2_STATE2_REG_1__SCAN_IN ? ~P2_PHYADDRPOINTER_REG_0__SCAN_IN : P2_STATE2_REG_0__SCAN_IN;
  assign new_n1398_ = (~P2_INSTADDRPOINTER_REG_1__SCAN_IN | ((new_n1374_ | ~P2_STATE2_REG_0__SCAN_IN) & ~new_n1376_ & (~new_n1375_ | ~P2_STATE2_REG_0__SCAN_IN))) & new_n1399_ & (~new_n1380_ | ~P2_REIP_REG_1__SCAN_IN);
  assign new_n1399_ = ~new_n1400_ & (~P2_EBX_REG_1__SCAN_IN | new_n1322_ | ~new_n1340_ | ~new_n1359_ | ~new_n1358_ | ~new_n1330_ | new_n1317_);
  assign new_n1400_ = P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign new_n1401_ = P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & (new_n1329_ | new_n1355_ | new_n1357_ | new_n1372_ | new_n1366_ | new_n1369_ | new_n1371_);
  assign new_n1402_ = new_n1403_ & (new_n1374_ | ~P2_STATE2_REG_0__SCAN_IN);
  assign new_n1403_ = (~new_n1330_ | ~new_n1377_ | ~new_n1350_ | ~new_n1356_ | new_n1322_ | ~new_n1340_) & ~new_n1404_ & (~new_n1330_ | ~new_n1377_ | ~new_n1350_ | ~new_n1356_ | ~new_n1340_ | new_n1378_);
  assign new_n1404_ = new_n1382_ & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n1405_ = (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | (~new_n1406_ & ~P2_STATE2_REG_3__SCAN_IN)) & (P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_2__SCAN_IN | (P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ^ (~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)));
  assign new_n1406_ = ~new_n1317_ & P2_STATE2_REG_0__SCAN_IN;
  assign new_n1407_ = P2_STATE2_REG_2__SCAN_IN & ~P2_STATE2_REG_0__SCAN_IN;
  assign new_n1408_ = ~new_n1314_ & new_n1405_ & (~new_n1407_ | (new_n1327_ & (new_n1383_ | (~new_n1386_ & ~new_n1387_))) | (~new_n1327_ & ~new_n1383_ & (new_n1386_ | new_n1387_)));
  assign new_n1409_ = (~P2_STATE2_REG_2__SCAN_IN | P2_STATE2_REG_0__SCAN_IN | (new_n1387_ & ~new_n1410_) | (~new_n1387_ & new_n1410_)) & (~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | (~P2_STATE2_REG_3__SCAN_IN & (new_n1317_ | ~P2_STATE2_REG_0__SCAN_IN))) & (~new_n1411_ | P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_2__SCAN_IN);
  assign new_n1410_ = (~new_n1384_ | (~new_n1373_ & P2_INSTADDRPOINTER_REG_2__SCAN_IN)) ^ (~new_n1385_ | (P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & (~new_n1328_ | ~new_n1365_)));
  assign new_n1411_ = P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ (P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  assign new_n1412_ = (~new_n1315_ | ~P2_INSTQUEUE_REG_0__1__SCAN_IN | (new_n1417_ & (~new_n1413_ | ~new_n1407_))) & (~new_n1414_ | ((~new_n1315_ | ~P2_INSTQUEUE_REG_0__1__SCAN_IN) & new_n1417_ & (~new_n1413_ | ~new_n1407_)));
  assign new_n1413_ = (~new_n1401_ & new_n1402_) ^ (new_n1398_ ^ (~new_n1390_ & (~new_n1328_ | ~new_n1388_) & (new_n1391_ | ~new_n1392_)));
  assign new_n1414_ = ~new_n1415_ & (~new_n1416_ | (new_n1407_ & (new_n1390_ | (new_n1328_ & new_n1388_) | (~new_n1391_ & new_n1392_)) & ((~new_n1390_ & (~new_n1328_ | ~new_n1388_)) | new_n1391_ | ~new_n1392_)));
  assign new_n1415_ = (~P2_INSTQUEUE_REG_0__0__SCAN_IN | ~new_n1316_ | new_n1322_) & new_n1316_ & ~P2_STATE2_REG_3__SCAN_IN & P2_STATE2_REG_2__SCAN_IN;
  assign new_n1416_ = (~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~new_n1406_ & ~P2_STATE2_REG_3__SCAN_IN)) & (P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_2__SCAN_IN);
  assign new_n1417_ = (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~new_n1406_ & ~P2_STATE2_REG_3__SCAN_IN)) & (new_n1418_ | P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_2__SCAN_IN);
  assign new_n1418_ = P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n1419_ = new_n1315_ & P2_INSTQUEUE_REG_0__5__SCAN_IN;
  assign new_n1420_ = (~new_n1315_ | ~P2_INSTQUEUE_REG_0__4__SCAN_IN) & (~new_n1406_ | ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  assign new_n1421_ = new_n1315_ & P2_INSTQUEUE_REG_0__2__SCAN_IN;
  assign new_n1422_ = new_n1315_ & ~new_n1423_;
  assign new_n1423_ = new_n1424_ & new_n1425_ & new_n1426_ & new_n1427_;
  assign new_n1424_ = (~P2_INSTQUEUE_REG_3__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_12__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_9__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1425_ = (~P2_INSTQUEUE_REG_4__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_11__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_1__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_15__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1426_ = (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUE_REG_13__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_7__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_14__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_8__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1427_ = (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_2__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_6__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_10__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_5__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1428_ = new_n1315_ & ~new_n1429_;
  assign new_n1429_ = new_n1430_ & new_n1434_ & new_n1435_ & (~P2_INSTQUEUE_REG_3__3__SCAN_IN | ~new_n1432_ | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_7__3__SCAN_IN | ~new_n1433_ | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1430_ = new_n1431_ & (~P2_INSTQUEUE_REG_0__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_9__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_1__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1431_ = (~P2_INSTQUEUE_REG_5__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_4__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_15__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_14__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1432_ = ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign new_n1433_ = P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign new_n1434_ = (~P2_INSTQUEUE_REG_8__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_6__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_10__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n1435_ = (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_2__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_12__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_13__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUE_REG_11__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1436_ = new_n1315_ & ~new_n1437_;
  assign new_n1437_ = new_n1438_ & new_n1440_ & new_n1441_ & (~P2_INSTQUEUE_REG_3__1__SCAN_IN | ~new_n1432_ | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_7__1__SCAN_IN | ~new_n1433_ | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1438_ = new_n1439_ & (~P2_INSTQUEUE_REG_1__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_15__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1439_ = (~P2_INSTQUEUE_REG_11__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_14__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_4__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_9__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1440_ = (~P2_INSTQUEUE_REG_5__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_2__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_12__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_13__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1441_ = (~P2_INSTQUEUE_REG_8__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_6__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_10__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n1442_ = new_n1315_ & P2_INSTQUEUE_REG_0__7__SCAN_IN;
  assign new_n1443_ = new_n1444_ & new_n1446_ & new_n1447_ & (~P2_INSTQUEUE_REG_3__0__SCAN_IN | ~new_n1432_ | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_7__0__SCAN_IN | ~new_n1433_ | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1444_ = new_n1445_ & (~P2_INSTQUEUE_REG_1__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_15__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1445_ = (~P2_INSTQUEUE_REG_11__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_14__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_4__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_9__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1446_ = (~P2_INSTQUEUE_REG_5__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_2__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_12__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_13__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1447_ = (~P2_INSTQUEUE_REG_8__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_6__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_10__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n1448_ = new_n1449_ & new_n1452_;
  assign new_n1449_ = new_n1450_ & new_n1451_ & (~P2_INSTQUEUE_REG_2__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_7__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1450_ = (~P2_INSTQUEUE_REG_11__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_6__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_8__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_10__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1451_ = (~P2_INSTQUEUE_REG_3__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_12__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_13__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1452_ = new_n1453_ & (~P2_INSTQUEUE_REG_0__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_9__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_1__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1453_ = (~P2_INSTQUEUE_REG_5__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_4__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_15__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_14__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1454_ = new_n1457_ & new_n1458_ & new_n1455_ & new_n1456_;
  assign new_n1455_ = (~P2_INSTQUEUE_REG_10__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_12__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_8__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_6__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1456_ = (~P2_INSTQUEUE_REG_3__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_7__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_2__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_5__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1457_ = (~P2_INSTQUEUE_REG_0__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_15__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_9__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_1__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1458_ = (~P2_INSTQUEUE_REG_14__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_13__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_4__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_11__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1459_ = new_n1315_ & ~new_n1460_;
  assign new_n1460_ = new_n1464_ & new_n1461_ & new_n1465_ & (~new_n1463_ | ~P2_INSTQUEUE_REG_1__7__SCAN_IN) & (~P2_INSTQUEUE_REG_11__7__SCAN_IN | ~new_n1432_ | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1461_ = new_n1462_ & (~P2_INSTQUEUE_REG_8__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_14__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_12__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1462_ = (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_10__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUE_REG_5__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_13__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_7__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1463_ = P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign new_n1464_ = (~P2_INSTQUEUE_REG_0__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_9__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_3__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_15__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1465_ = (~P2_INSTQUEUE_REG_4__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_2__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_6__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1466_ = new_n1316_ & (~new_n1467_ | ~new_n1469_ | ~new_n1470_ | (P2_INSTQUEUE_REG_4__0__SCAN_IN & new_n1432_ & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (P2_INSTQUEUE_REG_12__0__SCAN_IN & new_n1432_ & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1467_ = new_n1468_ & (~P2_INSTQUEUE_REG_2__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_13__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1468_ = (~P2_INSTQUEUE_REG_5__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_14__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_6__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_8__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1469_ = (~P2_INSTQUEUE_REG_10__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_3__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_1__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_15__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1470_ = (~P2_INSTQUEUE_REG_11__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_9__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_7__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n1471_ = new_n1474_ & new_n1472_ & new_n1475_ & (~new_n1463_ | ~P2_INSTQUEUE_REG_1__6__SCAN_IN) & (~P2_INSTQUEUE_REG_11__6__SCAN_IN | ~new_n1432_ | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1472_ = new_n1473_ & (~P2_INSTQUEUE_REG_8__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_14__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_12__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1473_ = (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_10__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUE_REG_5__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_13__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_7__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1474_ = (~P2_INSTQUEUE_REG_0__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_9__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_3__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_15__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1475_ = (~P2_INSTQUEUE_REG_4__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_2__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_6__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1476_ = new_n1477_ & new_n1479_ & new_n1480_ & (~P2_INSTQUEUE_REG_4__1__SCAN_IN | ~new_n1432_ | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_12__1__SCAN_IN | ~new_n1432_ | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1477_ = new_n1478_ & (~P2_INSTQUEUE_REG_2__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_6__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_0__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1478_ = (~P2_INSTQUEUE_REG_15__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_10__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_13__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_8__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1479_ = (~P2_INSTQUEUE_REG_1__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_3__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_14__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_5__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1480_ = (~P2_INSTQUEUE_REG_11__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_9__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_7__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n1481_ = new_n1316_ & (~new_n1482_ | ~new_n1484_ | ~new_n1485_ | (P2_INSTQUEUE_REG_4__2__SCAN_IN & new_n1432_ & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (P2_INSTQUEUE_REG_12__2__SCAN_IN & new_n1432_ & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1482_ = new_n1483_ & (~P2_INSTQUEUE_REG_2__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_13__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1483_ = (~P2_INSTQUEUE_REG_5__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_14__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_6__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_8__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1484_ = (~P2_INSTQUEUE_REG_10__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_3__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_1__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_15__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1485_ = (~P2_INSTQUEUE_REG_11__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_9__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_7__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n1486_ = new_n1316_ & (~new_n1489_ | ~new_n1490_ | ~new_n1487_ | ~new_n1488_);
  assign new_n1487_ = (~P2_INSTQUEUE_REG_9__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_7__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_14__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_11__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1488_ = (~P2_INSTQUEUE_REG_4__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_12__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_10__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_3__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1489_ = (~P2_INSTQUEUE_REG_13__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_6__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_2__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1490_ = (~P2_INSTQUEUE_REG_1__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_15__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_5__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_8__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1491_ = new_n1492_ & new_n1495_;
  assign new_n1492_ = new_n1493_ & new_n1494_ & (~P2_INSTQUEUE_REG_13__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_10__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1493_ = (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_3__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_7__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_15__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_9__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1494_ = (~P2_INSTQUEUE_REG_12__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_5__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_11__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1495_ = new_n1496_ & (~P2_INSTQUEUE_REG_6__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_14__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_4__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1496_ = (~P2_INSTQUEUE_REG_8__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_1__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_2__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1497_ = ~new_n1498_ & ~new_n1504_;
  assign new_n1498_ = new_n1502_ & new_n1499_ & new_n1503_;
  assign new_n1499_ = new_n1500_ & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_15__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_9__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_3__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1500_ = (new_n1501_ | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_5__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_11__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_7__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1501_ = P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_14__7__SCAN_IN : ~P2_INSTQUEUE_REG_6__7__SCAN_IN;
  assign new_n1502_ = (~P2_INSTQUEUE_REG_2__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_12__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_4__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1503_ = (~P2_INSTQUEUE_REG_13__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_10__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_1__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_8__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1504_ = new_n1505_ & new_n1508_ & ((~P2_INSTQUEUE_REG_3__0__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_11__0__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1505_ = new_n1507_ & new_n1506_ & ((~P2_INSTQUEUE_REG_0__0__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_8__0__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1506_ = ((~P2_INSTQUEUE_REG_1__0__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_9__0__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN)) & ((~P2_INSTQUEUE_REG_2__0__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_10__0__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1507_ = ((~P2_INSTQUEUE_REG_6__0__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_14__0__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_5__0__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_13__0__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1508_ = ((~P2_INSTQUEUE_REG_7__0__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_15__0__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_4__0__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_12__0__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1509_ = new_n1316_ & (~new_n1498_ | ~new_n1504_) & (new_n1322_ | new_n1498_ | new_n1504_);
  assign new_n1510_ = new_n1316_ & (~new_n1511_ | ~new_n1512_ | ~new_n1513_ | ~new_n1514_);
  assign new_n1511_ = (~P2_INSTQUEUE_REG_1__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_8__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_10__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_12__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1512_ = (~P2_INSTQUEUE_REG_13__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_2__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_4__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1513_ = (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_7__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_14__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_3__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_6__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1514_ = (~P2_INSTQUEUE_REG_15__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_9__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_11__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_5__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1515_ = new_n1516_ & new_n1519_ & ((~P2_INSTQUEUE_REG_3__1__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_11__1__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1516_ = new_n1518_ & new_n1517_ & ((~P2_INSTQUEUE_REG_0__1__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_8__1__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1517_ = ((~P2_INSTQUEUE_REG_1__1__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_9__1__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN)) & ((~P2_INSTQUEUE_REG_2__1__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_10__1__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1518_ = ((~P2_INSTQUEUE_REG_6__1__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_14__1__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_5__1__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_13__1__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1519_ = ((~P2_INSTQUEUE_REG_7__1__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_15__1__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_4__1__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_12__1__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1520_ = new_n1521_ & new_n1524_;
  assign new_n1521_ = new_n1522_ & new_n1523_ & (~P2_INSTQUEUE_REG_13__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_10__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1522_ = (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_3__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_7__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_14__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_9__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1523_ = (~P2_INSTQUEUE_REG_6__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_5__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_11__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1524_ = new_n1525_ & (~P2_INSTQUEUE_REG_12__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_15__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_4__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1525_ = (~P2_INSTQUEUE_REG_8__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_1__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_2__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1526_ = ~new_n1629_ ^ (~new_n1628_ & new_n1527_ & ~new_n1627_);
  assign new_n1527_ = new_n1528_ & ~new_n1626_;
  assign new_n1528_ = new_n1529_ & ~new_n1625_;
  assign new_n1529_ = new_n1530_ & ((~new_n1545_ & P2_INSTADDRPOINTER_REG_20__SCAN_IN) | (new_n1544_ & P2_EAX_REG_20__SCAN_IN) | (new_n1542_ & P2_REIP_REG_20__SCAN_IN));
  assign new_n1530_ = ~new_n1624_ & ~new_n1623_ & ~new_n1622_ & ~new_n1621_ & ~new_n1620_ & ~new_n1619_ & new_n1531_ & ~new_n1618_;
  assign new_n1531_ = ~new_n1617_ & ~new_n1616_ & ~new_n1615_ & ~new_n1614_ & ~new_n1613_ & (new_n1532_ | (~new_n1547_ & ~new_n1548_));
  assign new_n1532_ = new_n1533_ & (~new_n1541_ | (~new_n1545_ & P2_INSTADDRPOINTER_REG_7__SCAN_IN));
  assign new_n1533_ = ~new_n1534_ & new_n1540_;
  assign new_n1534_ = new_n1537_ & new_n1538_ & new_n1535_ & new_n1539_;
  assign new_n1535_ = (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUE_REG_12__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_11__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUE_REG_4__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (new_n1536_ | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1536_ = P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_13__7__SCAN_IN : ~P2_INSTQUEUE_REG_5__7__SCAN_IN;
  assign new_n1537_ = (~P2_INSTQUEUE_REG_1__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_10__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_8__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1538_ = (~P2_INSTQUEUE_REG_7__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_9__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_3__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1539_ = (~P2_INSTQUEUE_REG_14__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUE_REG_2__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_6__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_15__7__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1540_ = new_n1322_ & ~new_n1330_ & ~P2_STATE2_REG_3__SCAN_IN;
  assign new_n1541_ = (~new_n1542_ | ~P2_REIP_REG_7__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_7__SCAN_IN);
  assign new_n1542_ = new_n1543_ & new_n1322_ & new_n1330_;
  assign new_n1543_ = (~new_n1338_ | ~new_n1339_ | ~new_n1336_ | ~new_n1337_) & ~new_n1378_ & ~P2_STATE2_REG_3__SCAN_IN;
  assign new_n1544_ = new_n1335_ & ~P2_STATE2_REG_3__SCAN_IN;
  assign new_n1545_ = (new_n1317_ | ~new_n1543_) & (~new_n1330_ | ~new_n1546_) & (~new_n1546_ | new_n1330_ | ~new_n1317_);
  assign new_n1546_ = ~P2_STATE2_REG_3__SCAN_IN & (~new_n1325_ | ~new_n1326_ | ~new_n1323_ | ~new_n1324_);
  assign new_n1547_ = ~new_n1533_ & new_n1541_ & (new_n1545_ | ~P2_INSTADDRPOINTER_REG_7__SCAN_IN);
  assign new_n1548_ = ~new_n1549_ & (new_n1557_ | (~new_n1558_ & (new_n1566_ | (~new_n1567_ & (new_n1575_ | new_n1576_)))));
  assign new_n1549_ = new_n1550_ & ((~new_n1545_ & P2_INSTADDRPOINTER_REG_6__SCAN_IN) | (new_n1544_ & P2_EAX_REG_6__SCAN_IN) | (new_n1542_ & P2_REIP_REG_6__SCAN_IN));
  assign new_n1550_ = ~new_n1551_ & new_n1322_ & ~new_n1330_ & ~P2_STATE2_REG_3__SCAN_IN;
  assign new_n1551_ = new_n1552_ & new_n1553_ & new_n1556_ & new_n1554_ & new_n1555_;
  assign new_n1552_ = (~P2_INSTQUEUE_REG_1__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_10__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_8__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1553_ = (~P2_INSTQUEUE_REG_7__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_9__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_3__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1554_ = (~P2_INSTQUEUE_REG_12__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_11__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1555_ = (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_13__6__SCAN_IN : ~P2_INSTQUEUE_REG_5__6__SCAN_IN)) & (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUE_REG_4__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1556_ = (~P2_INSTQUEUE_REG_14__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUE_REG_2__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_6__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_15__6__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1557_ = ~new_n1550_ & (new_n1545_ | ~P2_INSTADDRPOINTER_REG_6__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_6__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_6__SCAN_IN);
  assign new_n1558_ = new_n1559_ & ((~new_n1545_ & P2_INSTADDRPOINTER_REG_5__SCAN_IN) | (new_n1544_ & P2_EAX_REG_5__SCAN_IN) | (new_n1542_ & P2_REIP_REG_5__SCAN_IN));
  assign new_n1559_ = ~new_n1560_ & new_n1322_ & ~new_n1330_ & ~P2_STATE2_REG_3__SCAN_IN;
  assign new_n1560_ = new_n1561_ & new_n1562_ & new_n1565_ & new_n1563_ & new_n1564_;
  assign new_n1561_ = (~P2_INSTQUEUE_REG_8__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_3__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1562_ = (~P2_INSTQUEUE_REG_4__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_1__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_10__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_12__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1563_ = (~P2_INSTQUEUE_REG_11__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ? ~P2_INSTQUEUE_REG_13__5__SCAN_IN : ~P2_INSTQUEUE_REG_5__5__SCAN_IN));
  assign new_n1564_ = (~P2_INSTQUEUE_REG_9__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_7__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1565_ = (~P2_INSTQUEUE_REG_14__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUE_REG_2__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_6__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_15__5__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1566_ = ~new_n1559_ & (new_n1545_ | ~P2_INSTADDRPOINTER_REG_5__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_5__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_5__SCAN_IN);
  assign new_n1567_ = new_n1568_ & ((~new_n1545_ & P2_INSTADDRPOINTER_REG_4__SCAN_IN) | (new_n1544_ & P2_EAX_REG_4__SCAN_IN) | (new_n1542_ & P2_REIP_REG_4__SCAN_IN));
  assign new_n1568_ = ~new_n1569_ & new_n1322_ & ~new_n1330_ & ~P2_STATE2_REG_3__SCAN_IN;
  assign new_n1569_ = new_n1573_ & new_n1574_ & new_n1570_ & new_n1571_ & new_n1572_;
  assign new_n1570_ = (~P2_INSTQUEUE_REG_14__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_12__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_10__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1571_ = (~P2_INSTQUEUE_REG_5__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_9__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUE_REG_4__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUE_REG_7__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1572_ = (~P2_INSTQUEUE_REG_13__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_2__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1573_ = (~P2_INSTQUEUE_REG_11__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__4__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_6__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1574_ = (~P2_INSTQUEUE_REG_8__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_15__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_3__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_1__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1575_ = ~new_n1568_ & (new_n1545_ | ~P2_INSTADDRPOINTER_REG_4__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_4__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_4__SCAN_IN);
  assign new_n1576_ = (new_n1604_ | ((new_n1595_ | ((new_n1586_ | new_n1577_ | new_n1579_) & (new_n1593_ | (new_n1586_ & (new_n1577_ | new_n1579_))))) & (new_n1602_ | (new_n1595_ & (new_n1586_ | new_n1577_ | new_n1579_) & (new_n1593_ | (new_n1586_ & (new_n1577_ | new_n1579_))))))) & (new_n1606_ | (new_n1604_ & (new_n1595_ | ((new_n1586_ | new_n1577_ | new_n1579_) & (new_n1593_ | (new_n1586_ & (new_n1577_ | new_n1579_))))) & (new_n1602_ | (new_n1595_ & (new_n1586_ | new_n1577_ | new_n1579_) & (new_n1593_ | (new_n1586_ & (new_n1577_ | new_n1579_)))))));
  assign new_n1577_ = (~P2_INSTADDRPOINTER_REG_0__SCAN_IN | ((new_n1317_ | ~new_n1543_) & (~new_n1330_ | ~new_n1546_) & (~new_n1546_ | new_n1330_ | ~new_n1317_))) & new_n1578_ & (~P2_REIP_REG_0__SCAN_IN | ~new_n1543_ | ~new_n1322_ | ~new_n1330_);
  assign new_n1578_ = ~P2_STATE2_REG_3__SCAN_IN & (~P2_EAX_REG_0__SCAN_IN | ~new_n1338_ | ~new_n1339_ | ~new_n1336_ | ~new_n1337_);
  assign new_n1579_ = (new_n1580_ | ~new_n1322_ | new_n1330_ | P2_STATE2_REG_3__SCAN_IN) & (new_n1330_ | ~new_n1317_ | new_n1322_ | P2_STATE2_REG_3__SCAN_IN) & (~P2_STATE2_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (~new_n1335_ | P2_STATE2_REG_3__SCAN_IN);
  assign new_n1580_ = new_n1584_ & new_n1585_ & new_n1581_ & new_n1582_ & new_n1583_;
  assign new_n1581_ = (~P2_INSTQUEUE_REG_4__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_3__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_13__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_12__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1582_ = (~P2_INSTQUEUE_REG_7__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_5__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_9__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n1583_ = (~P2_INSTQUEUE_REG_2__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_6__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1584_ = (~P2_INSTQUEUE_REG_14__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_8__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_11__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1585_ = (~P2_INSTQUEUE_REG_0__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_1__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_10__0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_15__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1586_ = (new_n1587_ | ~new_n1322_ | new_n1330_ | P2_STATE2_REG_3__SCAN_IN) & (~new_n1543_ | (~new_n1330_ & new_n1317_)) & (~P2_STATE2_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~new_n1330_ | new_n1322_ | P2_STATE2_REG_3__SCAN_IN);
  assign new_n1587_ = new_n1591_ & new_n1592_ & new_n1588_ & new_n1589_ & new_n1590_;
  assign new_n1588_ = (~P2_INSTQUEUE_REG_4__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_15__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_2__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_1__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1589_ = (~P2_INSTQUEUE_REG_7__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_5__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_9__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n1590_ = (~P2_INSTQUEUE_REG_13__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_8__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1591_ = (~P2_INSTQUEUE_REG_3__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_11__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_10__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1592_ = (~P2_INSTQUEUE_REG_14__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_12__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_0__1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_6__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1593_ = (~P2_INSTADDRPOINTER_REG_1__SCAN_IN | ((new_n1317_ | ~new_n1543_) & (new_n1330_ | ~new_n1317_ | new_n1322_ | P2_STATE2_REG_3__SCAN_IN) & (~new_n1330_ | new_n1322_ | P2_STATE2_REG_3__SCAN_IN))) & ~new_n1594_ & (~P2_REIP_REG_1__SCAN_IN | ~new_n1543_ | ~new_n1322_ | ~new_n1330_);
  assign new_n1594_ = P2_EAX_REG_1__SCAN_IN & ~P2_STATE2_REG_3__SCAN_IN & new_n1338_ & new_n1339_ & new_n1336_ & new_n1337_;
  assign new_n1595_ = (new_n1596_ | ~new_n1322_ | new_n1330_ | P2_STATE2_REG_3__SCAN_IN) & (~P2_STATE2_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (new_n1330_ | ~new_n1317_ | new_n1322_ | P2_STATE2_REG_3__SCAN_IN);
  assign new_n1596_ = new_n1600_ & new_n1601_ & new_n1597_ & new_n1598_ & new_n1599_;
  assign new_n1597_ = (~P2_INSTQUEUE_REG_5__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_1__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_7__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1598_ = (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUE_REG_12__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_13__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_3__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUE_REG_9__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1599_ = (~P2_INSTQUEUE_REG_2__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_14__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1600_ = (~P2_INSTQUEUE_REG_11__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_8__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1601_ = (~P2_INSTQUEUE_REG_10__2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_15__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_6__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_4__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1602_ = (~P2_INSTADDRPOINTER_REG_2__SCAN_IN | ((new_n1317_ | ~new_n1543_) & (new_n1330_ | ~new_n1317_ | new_n1322_ | P2_STATE2_REG_3__SCAN_IN) & (~new_n1330_ | new_n1322_ | P2_STATE2_REG_3__SCAN_IN))) & ~new_n1603_ & (~P2_REIP_REG_2__SCAN_IN | ~new_n1543_ | ~new_n1322_ | ~new_n1330_);
  assign new_n1603_ = P2_EAX_REG_2__SCAN_IN & ~P2_STATE2_REG_3__SCAN_IN & new_n1338_ & new_n1339_ & new_n1336_ & new_n1337_;
  assign new_n1604_ = (~P2_INSTADDRPOINTER_REG_3__SCAN_IN | ((new_n1317_ | ~new_n1543_) & (new_n1330_ | ~new_n1317_ | new_n1322_ | P2_STATE2_REG_3__SCAN_IN) & (~new_n1330_ | new_n1322_ | P2_STATE2_REG_3__SCAN_IN))) & ~new_n1605_ & (~P2_REIP_REG_3__SCAN_IN | ~new_n1543_ | ~new_n1322_ | ~new_n1330_);
  assign new_n1605_ = P2_EAX_REG_3__SCAN_IN & ~P2_STATE2_REG_3__SCAN_IN & new_n1338_ & new_n1339_ & new_n1336_ & new_n1337_;
  assign new_n1606_ = (~P2_STATE2_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) & (new_n1607_ | ~new_n1322_ | new_n1330_ | P2_STATE2_REG_3__SCAN_IN);
  assign new_n1607_ = new_n1611_ & new_n1612_ & new_n1608_ & new_n1609_ & new_n1610_;
  assign new_n1608_ = (~P2_INSTQUEUE_REG_12__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_7__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUE_REG_3__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUE_REG_10__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n1609_ = (~P2_INSTQUEUE_REG_13__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_5__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P2_INSTQUEUE_REG_9__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n1610_ = (~P2_INSTQUEUE_REG_2__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_15__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1611_ = (~P2_INSTQUEUE_REG_11__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_0__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_6__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n1612_ = (~P2_INSTQUEUE_REG_8__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUE_REG_4__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_14__3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUE_REG_1__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n1613_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_8__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_8__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_8__SCAN_IN) & (~new_n1540_ | new_n1443_);
  assign new_n1614_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_9__SCAN_IN) & (~new_n1540_ | new_n1437_) & (~new_n1544_ | ~P2_EAX_REG_9__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_9__SCAN_IN);
  assign new_n1615_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_10__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_10__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_10__SCAN_IN) & (~new_n1540_ | new_n1448_);
  assign new_n1616_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_11__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_11__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_11__SCAN_IN) & (~new_n1540_ | new_n1429_);
  assign new_n1617_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_12__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_12__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_12__SCAN_IN) & (~new_n1540_ | new_n1454_);
  assign new_n1618_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_13__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_13__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_13__SCAN_IN) & (~new_n1540_ | new_n1423_);
  assign new_n1619_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_14__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_14__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_14__SCAN_IN) & (~new_n1540_ | new_n1471_);
  assign new_n1620_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_15__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_15__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_15__SCAN_IN) & (~new_n1540_ | new_n1460_);
  assign new_n1621_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_16__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_16__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_16__SCAN_IN);
  assign new_n1622_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_17__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_17__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_17__SCAN_IN);
  assign new_n1623_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_18__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_18__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_18__SCAN_IN);
  assign new_n1624_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_19__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_19__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_19__SCAN_IN);
  assign new_n1625_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_21__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_21__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_21__SCAN_IN);
  assign new_n1626_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_22__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_22__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_22__SCAN_IN);
  assign new_n1627_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_23__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_23__SCAN_IN);
  assign new_n1628_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_24__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_24__SCAN_IN);
  assign new_n1629_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_25__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_25__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_25__SCAN_IN);
  assign new_n1630_ = (new_n1632_ | ~new_n1316_ | ~new_n1322_) & ((~new_n1631_ & new_n1632_) | ~new_n1316_ | new_n1322_ | (new_n1631_ & ~new_n1632_));
  assign new_n1631_ = new_n1497_ & ~new_n1515_;
  assign new_n1632_ = new_n1633_ & new_n1636_ & ((~P2_INSTQUEUE_REG_3__2__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_11__2__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1633_ = new_n1635_ & new_n1634_ & ((~P2_INSTQUEUE_REG_0__2__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_8__2__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1634_ = ((~P2_INSTQUEUE_REG_1__2__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_9__2__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN)) & ((~P2_INSTQUEUE_REG_2__2__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_10__2__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1635_ = ((~P2_INSTQUEUE_REG_6__2__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_14__2__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_5__2__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_13__2__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1636_ = ((~P2_INSTQUEUE_REG_7__2__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_15__2__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_4__2__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_12__2__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1637_ = ~new_n1638_ & (new_n1640_ | ((~new_n1700_ | (new_n1699_ & new_n1486_) | (~new_n1699_ & ~new_n1486_)) & ((~new_n1700_ & (~new_n1699_ ^ new_n1486_)) | (~new_n1641_ & (new_n1647_ | ~new_n1698_)))));
  assign new_n1638_ = new_n1639_ & (~new_n1309_ | new_n1520_) & (new_n1309_ | (new_n1316_ & ~new_n1520_));
  assign new_n1639_ = new_n1529_ ^ ~new_n1625_;
  assign new_n1640_ = ~new_n1639_ & (new_n1309_ ? ~new_n1520_ : (~new_n1316_ | new_n1520_));
  assign new_n1641_ = new_n1646_ & (new_n1624_ | new_n1623_ | ~new_n1642_ | new_n1622_) & (~new_n1624_ | (~new_n1623_ & new_n1642_ & ~new_n1622_));
  assign new_n1642_ = new_n1643_ & ~new_n1621_;
  assign new_n1643_ = new_n1644_ & ~new_n1620_;
  assign new_n1644_ = new_n1645_ & ~new_n1619_;
  assign new_n1645_ = new_n1531_ & ~new_n1618_;
  assign new_n1646_ = (new_n1481_ & ~new_n1476_ & new_n1466_ & new_n1459_ & new_n1311_ & ~new_n1471_) ? new_n1491_ : (new_n1316_ & ~new_n1491_);
  assign new_n1647_ = new_n1691_ & (new_n1695_ | (~new_n1648_ & ~new_n1696_) | ((~new_n1687_ | (new_n1649_ & ~new_n1697_)) & ~new_n1690_ & (~new_n1648_ | ~new_n1696_)));
  assign new_n1648_ = new_n1643_ ^ ~new_n1621_;
  assign new_n1649_ = (~new_n1650_ | ~new_n1686_) & ((~new_n1650_ & ~new_n1686_) | new_n1652_ | (new_n1685_ & (new_n1655_ | ~new_n1682_)));
  assign new_n1650_ = new_n1422_ ^ (~new_n1454_ & new_n1651_ & new_n1428_);
  assign new_n1651_ = ~new_n1448_ & new_n1436_ & ~new_n1443_ & new_n1312_ & new_n1442_;
  assign new_n1652_ = (new_n1653_ ^ new_n1617_) & ((new_n1651_ & ~new_n1429_ & new_n1316_ & ~new_n1322_) ? ~new_n1454_ : (new_n1454_ | ~new_n1316_ | new_n1322_));
  assign new_n1653_ = new_n1654_ & ~new_n1616_;
  assign new_n1654_ = ~new_n1615_ & ~new_n1614_ & ~new_n1613_ & (new_n1532_ | (~new_n1547_ & ~new_n1548_));
  assign new_n1655_ = ~new_n1656_ & ((~new_n1658_ & ~new_n1681_) | ((~new_n1658_ | ~new_n1681_) & (new_n1659_ | (new_n1680_ & (~new_n1677_ | (~new_n1661_ & new_n1675_))))));
  assign new_n1656_ = new_n1657_ & (new_n1448_ | ~new_n1315_ | new_n1437_ | new_n1443_ | ~new_n1312_ | ~P2_INSTQUEUE_REG_0__7__SCAN_IN) & ((new_n1315_ & ~new_n1437_ & ~new_n1443_ & new_n1312_ & P2_INSTQUEUE_REG_0__7__SCAN_IN) | (new_n1315_ & ~new_n1448_));
  assign new_n1657_ = ~new_n1615_ ^ (~new_n1614_ & ~new_n1613_ & (new_n1532_ | (~new_n1547_ & ~new_n1548_)));
  assign new_n1658_ = new_n1436_ ^ (~new_n1443_ & new_n1312_ & new_n1442_);
  assign new_n1659_ = ~new_n1660_ & ((new_n1312_ & new_n1315_ & P2_INSTQUEUE_REG_0__7__SCAN_IN) ? ~new_n1443_ : (~new_n1315_ | new_n1443_));
  assign new_n1660_ = ~new_n1613_ ^ (new_n1532_ | (~new_n1547_ & ~new_n1548_));
  assign new_n1661_ = (new_n1672_ | (new_n1419_ ^ (~new_n1662_ & ~new_n1420_))) & (new_n1673_ | (new_n1662_ ^ new_n1420_)) & ((new_n1673_ & (~new_n1662_ | ~new_n1420_) & (new_n1662_ | new_n1420_)) | ((new_n1663_ | new_n1674_) & (~new_n1665_ | (new_n1663_ & new_n1674_))));
  assign new_n1662_ = ~new_n1313_ & (new_n1408_ | (new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_)));
  assign new_n1663_ = new_n1664_ ^ ((~new_n1412_ | (~new_n1409_ & new_n1421_)) & (~new_n1409_ | new_n1421_));
  assign new_n1664_ = new_n1314_ ^ (~new_n1405_ | (new_n1407_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_))));
  assign new_n1665_ = (~new_n1667_ | ((new_n1412_ ^ (~new_n1409_ ^ new_n1421_)) & (~new_n1669_ | ~new_n1670_ | ~new_n1671_) & (~new_n1666_ | (~new_n1669_ & (~new_n1670_ | ~new_n1671_))))) & ((~new_n1412_ & (new_n1409_ | ~new_n1421_) & (~new_n1409_ | new_n1421_)) | (new_n1412_ & (new_n1409_ ^ new_n1421_)) | ((~new_n1669_ | ~new_n1670_ | ~new_n1671_) & (~new_n1666_ | (~new_n1669_ & (~new_n1670_ | ~new_n1671_)))));
  assign new_n1666_ = ~new_n1414_ ^ ((~new_n1315_ | ~P2_INSTQUEUE_REG_0__1__SCAN_IN) ^ (~new_n1417_ | (new_n1413_ & new_n1407_)));
  assign new_n1667_ = new_n1602_ ^ (new_n1595_ ^ ((new_n1668_ & ~new_n1586_) | (~new_n1593_ & (new_n1668_ | ~new_n1586_))));
  assign new_n1668_ = ~new_n1577_ & ~new_n1579_;
  assign new_n1669_ = new_n1593_ ^ (~new_n1668_ ^ ~new_n1586_);
  assign new_n1670_ = ~new_n1415_ ^ (~new_n1416_ | (new_n1407_ & (new_n1390_ | (new_n1328_ & new_n1388_) | (~new_n1391_ & new_n1392_)) & ((~new_n1390_ & (~new_n1328_ | ~new_n1388_)) | new_n1391_ | ~new_n1392_)));
  assign new_n1671_ = new_n1577_ ^ new_n1579_;
  assign new_n1672_ = (new_n1567_ | (~new_n1575_ & ~new_n1576_)) ^ (~new_n1558_ & ~new_n1566_);
  assign new_n1673_ = ~new_n1576_ ^ (~new_n1567_ & ~new_n1575_);
  assign new_n1674_ = new_n1606_ ^ (new_n1604_ ^ ((~new_n1595_ & ((new_n1668_ & ~new_n1586_) | (~new_n1593_ & (new_n1668_ | ~new_n1586_)))) | (~new_n1602_ & (~new_n1595_ | (new_n1668_ & ~new_n1586_) | (~new_n1593_ & (new_n1668_ | ~new_n1586_))))));
  assign new_n1675_ = (~new_n1672_ | (~new_n1662_ & ~new_n1420_ & P2_INSTQUEUE_REG_0__5__SCAN_IN & new_n1316_ & ~new_n1322_) | ((new_n1662_ | new_n1420_) & (~P2_INSTQUEUE_REG_0__5__SCAN_IN | ~new_n1316_ | new_n1322_))) & (~new_n1676_ | (P2_INSTQUEUE_REG_0__6__SCAN_IN & ~new_n1662_ & ~new_n1420_ & P2_INSTQUEUE_REG_0__5__SCAN_IN & new_n1316_ & ~new_n1322_) | ((new_n1662_ | new_n1420_ | ~P2_INSTQUEUE_REG_0__5__SCAN_IN | ~new_n1316_ | new_n1322_) & (~P2_INSTQUEUE_REG_0__6__SCAN_IN | ~new_n1316_ | new_n1322_)));
  assign new_n1676_ = (~new_n1549_ & ~new_n1557_) ^ (new_n1558_ | (~new_n1566_ & (new_n1567_ | (~new_n1575_ & ~new_n1576_))));
  assign new_n1677_ = (new_n1678_ | ((new_n1315_ & P2_INSTQUEUE_REG_0__7__SCAN_IN) ^ (P2_INSTQUEUE_REG_0__6__SCAN_IN & new_n1315_ & P2_INSTQUEUE_REG_0__5__SCAN_IN & ~new_n1662_ & ~new_n1420_))) & (new_n1676_ | ((new_n1315_ & P2_INSTQUEUE_REG_0__5__SCAN_IN & ~new_n1662_ & ~new_n1420_) ? ~P2_INSTQUEUE_REG_0__6__SCAN_IN : (new_n1315_ & P2_INSTQUEUE_REG_0__6__SCAN_IN)));
  assign new_n1678_ = new_n1679_ ^ (new_n1549_ | (~new_n1557_ & (new_n1558_ | (~new_n1566_ & (new_n1567_ | (~new_n1575_ & ~new_n1576_))))));
  assign new_n1679_ = (~new_n1534_ & new_n1540_) ^ ((~new_n1545_ & P2_INSTADDRPOINTER_REG_7__SCAN_IN) | (new_n1544_ & P2_EAX_REG_7__SCAN_IN) | (new_n1542_ & P2_REIP_REG_7__SCAN_IN));
  assign new_n1680_ = (~new_n1660_ | (~new_n1443_ & new_n1312_ & new_n1315_ & P2_INSTQUEUE_REG_0__7__SCAN_IN) | ((~new_n1315_ | new_n1443_) & (~new_n1312_ | ~new_n1315_ | ~P2_INSTQUEUE_REG_0__7__SCAN_IN))) & (~new_n1678_ | (new_n1312_ & new_n1315_ & P2_INSTQUEUE_REG_0__7__SCAN_IN) | (~new_n1312_ & (~new_n1315_ | ~P2_INSTQUEUE_REG_0__7__SCAN_IN)));
  assign new_n1681_ = ~new_n1614_ ^ (~new_n1613_ & (new_n1532_ | (~new_n1547_ & ~new_n1548_)));
  assign new_n1682_ = ~new_n1683_ & (new_n1684_ | (new_n1651_ ^ new_n1428_));
  assign new_n1683_ = ~new_n1657_ & ((new_n1315_ & ~new_n1437_ & ~new_n1443_ & new_n1312_ & P2_INSTQUEUE_REG_0__7__SCAN_IN) ? ~new_n1448_ : (~new_n1315_ | new_n1448_));
  assign new_n1684_ = new_n1654_ ^ ~new_n1616_;
  assign new_n1685_ = (~new_n1684_ | (new_n1651_ & ~new_n1429_ & new_n1316_ & ~new_n1322_) | (~new_n1651_ & (new_n1429_ | ~new_n1316_ | new_n1322_))) & ((new_n1653_ & ~new_n1617_) | (~new_n1653_ & new_n1617_) | (~new_n1454_ & new_n1651_ & ~new_n1429_ & new_n1316_ & ~new_n1322_) | ((new_n1454_ | ~new_n1316_ | new_n1322_) & (~new_n1651_ | new_n1429_ | ~new_n1316_ | new_n1322_)));
  assign new_n1686_ = new_n1531_ ^ ~new_n1618_;
  assign new_n1687_ = (new_n1689_ | (new_n1311_ ? new_n1471_ : (new_n1315_ & ~new_n1471_))) & (new_n1688_ | ((new_n1311_ & ~new_n1471_) ^ (new_n1315_ & ~new_n1460_)));
  assign new_n1688_ = new_n1644_ ^ ~new_n1620_;
  assign new_n1689_ = new_n1645_ ^ ~new_n1619_;
  assign new_n1690_ = new_n1688_ & (~new_n1459_ | ~new_n1311_ | new_n1471_) & (new_n1459_ | (new_n1311_ & ~new_n1471_));
  assign new_n1691_ = ~new_n1692_ & (~new_n1694_ | (new_n1310_ & new_n1481_) | (~new_n1310_ & ~new_n1481_));
  assign new_n1692_ = new_n1693_ & (new_n1476_ | ~new_n1466_ | ~new_n1459_ | ~new_n1311_ | new_n1471_) & ((new_n1316_ & ~new_n1476_) | (new_n1466_ & new_n1459_ & new_n1311_ & ~new_n1471_));
  assign new_n1693_ = ~new_n1622_ ^ (~new_n1621_ & ~new_n1620_ & new_n1645_ & ~new_n1619_);
  assign new_n1694_ = ~new_n1623_ ^ (~new_n1622_ & ~new_n1621_ & ~new_n1620_ & new_n1645_ & ~new_n1619_);
  assign new_n1695_ = ~new_n1693_ & ((new_n1466_ & new_n1459_ & new_n1311_ & ~new_n1471_) ? ~new_n1476_ : (~new_n1316_ | new_n1476_));
  assign new_n1696_ = new_n1466_ ^ (new_n1459_ & new_n1311_ & ~new_n1471_);
  assign new_n1697_ = new_n1689_ & (~new_n1311_ | new_n1471_) & (new_n1311_ | (new_n1315_ & ~new_n1471_));
  assign new_n1698_ = (new_n1646_ | (~new_n1624_ ^ (~new_n1623_ & new_n1642_ & ~new_n1622_))) & ((~new_n1623_ ^ (new_n1642_ & ~new_n1622_)) | (~new_n1310_ ^ ~new_n1481_));
  assign new_n1699_ = ~new_n1491_ & new_n1310_ & new_n1481_;
  assign new_n1700_ = new_n1530_ ^ ((~new_n1545_ & P2_INSTADDRPOINTER_REG_20__SCAN_IN) | (new_n1544_ & P2_EAX_REG_20__SCAN_IN) | (new_n1542_ & P2_REIP_REG_20__SCAN_IN));
  assign new_n1701_ = ~new_n1628_ ^ (new_n1527_ & ~new_n1627_);
  assign new_n1702_ = ~new_n1704_ ^ (new_n1509_ & (new_n1703_ | (new_n1510_ & new_n1309_ & ~new_n1520_)));
  assign new_n1703_ = new_n1497_ & new_n1316_ & new_n1322_;
  assign new_n1704_ = (new_n1515_ | ~new_n1316_ | ~new_n1322_) & ((~new_n1497_ & new_n1515_) | ~new_n1316_ | new_n1322_ | (new_n1497_ & ~new_n1515_));
  assign new_n1705_ = new_n1527_ ^ ~new_n1627_;
  assign new_n1706_ = ~new_n1707_ ^ (new_n1510_ & new_n1309_ & ~new_n1520_);
  assign new_n1707_ = ~new_n1703_ & new_n1509_;
  assign new_n1708_ = new_n1709_ & (~new_n1510_ | ~new_n1309_ | new_n1520_) & (new_n1510_ | (new_n1309_ & ~new_n1520_));
  assign new_n1709_ = new_n1528_ ^ ~new_n1626_;
  assign new_n1710_ = ~new_n1709_ & (~new_n1510_ ^ (new_n1309_ & ~new_n1520_));
  assign new_n1711_ = ~new_n1712_ & (~new_n1720_ | (~new_n1726_ & new_n1727_) | (new_n1726_ & ~new_n1727_));
  assign new_n1712_ = new_n1713_ & (((new_n1308_ | ((new_n1632_ | ~new_n1316_ | ~new_n1322_) & ((~new_n1631_ & new_n1632_) | (new_n1631_ & ~new_n1632_) | ~new_n1316_ | new_n1322_))) & (new_n1632_ | ~new_n1316_ | ~new_n1322_ | new_n1631_ | new_n1322_)) | ((new_n1715_ | ~new_n1316_ | ~new_n1322_) & (~new_n1316_ | new_n1322_ | (~new_n1715_ & new_n1631_ & ~new_n1632_) | (new_n1715_ & (~new_n1631_ | new_n1632_))))) & ((~new_n1308_ & ((~new_n1632_ & new_n1316_ & new_n1322_) | ((new_n1631_ | ~new_n1632_) & (~new_n1631_ | new_n1632_) & new_n1316_ & ~new_n1322_))) | (~new_n1632_ & new_n1316_ & new_n1322_ & ~new_n1631_ & ~new_n1322_) | (~new_n1715_ & new_n1316_ & new_n1322_) | (new_n1316_ & ~new_n1322_ & (new_n1715_ | ~new_n1631_ | new_n1632_) & (~new_n1715_ | (new_n1631_ & ~new_n1632_))));
  assign new_n1713_ = ~new_n1714_ ^ (~new_n1629_ & ~new_n1628_ & new_n1527_ & ~new_n1627_);
  assign new_n1714_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_26__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_26__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_26__SCAN_IN);
  assign new_n1715_ = new_n1716_ & new_n1719_ & ((~P2_INSTQUEUE_REG_3__3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_11__3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1716_ = new_n1718_ & new_n1717_ & ((~P2_INSTQUEUE_REG_0__3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_8__3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1717_ = ((~P2_INSTQUEUE_REG_1__3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_9__3__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN)) & ((~P2_INSTQUEUE_REG_2__3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_10__3__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1718_ = ((~P2_INSTQUEUE_REG_6__3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_14__3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_5__3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_13__3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1719_ = ((~P2_INSTQUEUE_REG_7__3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_15__3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_4__3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_12__3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1720_ = ((((~new_n1308_ & ((~new_n1632_ & new_n1316_ & new_n1322_) | ((new_n1631_ | ~new_n1632_) & new_n1316_ & ~new_n1322_ & (~new_n1631_ | new_n1632_)))) | (~new_n1632_ & new_n1316_ & new_n1322_ & ~new_n1631_ & ~new_n1322_)) & ((~new_n1715_ & new_n1316_ & new_n1322_) | (new_n1316_ & ~new_n1322_ & (new_n1715_ | ~new_n1631_ | new_n1632_) & (~new_n1715_ | (new_n1631_ & ~new_n1632_))))) | (new_n1316_ & ~new_n1322_ & (~new_n1631_ | new_n1632_) & ~new_n1715_ & new_n1322_)) ^ ((~new_n1721_ & new_n1316_ & new_n1322_) | (new_n1316_ & ~new_n1322_ & (new_n1721_ | new_n1715_ | ~new_n1631_ | new_n1632_) & (~new_n1721_ | (~new_n1715_ & new_n1631_ & ~new_n1632_))));
  assign new_n1721_ = new_n1722_ & new_n1725_ & ((~P2_INSTQUEUE_REG_3__4__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_11__4__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1722_ = new_n1724_ & new_n1723_ & ((~P2_INSTQUEUE_REG_0__4__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_8__4__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1723_ = ((~P2_INSTQUEUE_REG_1__4__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_9__4__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN)) & ((~P2_INSTQUEUE_REG_2__4__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_10__4__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1724_ = ((~P2_INSTQUEUE_REG_6__4__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_14__4__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_5__4__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_13__4__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1725_ = ((~P2_INSTQUEUE_REG_7__4__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_15__4__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_4__4__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_12__4__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1726_ = ~new_n1714_ & ~new_n1629_ & ~new_n1628_ & new_n1527_ & ~new_n1627_;
  assign new_n1727_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_27__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_27__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_27__SCAN_IN);
  assign new_n1728_ = ~new_n1713_ & (((new_n1308_ | ((new_n1632_ | ~new_n1316_ | ~new_n1322_) & ((~new_n1631_ & new_n1632_) | (new_n1631_ & ~new_n1632_) | ~new_n1316_ | new_n1322_))) & (new_n1632_ | ~new_n1316_ | ~new_n1322_ | new_n1631_ | new_n1322_)) ^ ((~new_n1715_ & new_n1316_ & new_n1322_) | (new_n1316_ & ~new_n1322_ & (new_n1715_ | ~new_n1631_ | new_n1632_) & (~new_n1715_ | (new_n1631_ & ~new_n1632_)))));
  assign new_n1729_ = (~new_n1730_ | ~new_n1743_) & (~new_n1747_ | (~new_n1731_ & new_n1748_) | (new_n1731_ & ~new_n1748_));
  assign new_n1730_ = (((~new_n1733_ & new_n1316_ & new_n1322_) ? ((new_n1732_ & ~new_n1738_) | ~new_n1316_ | new_n1322_) : ((~new_n1733_ | (new_n1732_ & ~new_n1738_)) & new_n1316_ & ~new_n1322_ & (new_n1733_ | ~new_n1732_ | new_n1738_))) | (~new_n1738_ & new_n1316_ & new_n1322_ & ~new_n1732_ & ~new_n1322_) | (~new_n1731_ & ((~new_n1738_ & new_n1316_ & new_n1322_) | ((new_n1732_ | ~new_n1738_) & (~new_n1732_ | new_n1738_) & new_n1316_ & ~new_n1322_)))) & ((~new_n1733_ & new_n1316_ & new_n1322_ & (~new_n1732_ | new_n1738_) & ~new_n1322_) | ((new_n1733_ | ~new_n1316_ | ~new_n1322_) & ((new_n1733_ & (~new_n1732_ | new_n1738_)) | ~new_n1316_ | new_n1322_ | (~new_n1733_ & new_n1732_ & ~new_n1738_))) | ((new_n1738_ | ~new_n1316_ | ~new_n1322_ | new_n1732_ | new_n1322_) & (new_n1731_ | ((new_n1738_ | ~new_n1316_ | ~new_n1322_) & ((~new_n1732_ & new_n1738_) | (new_n1732_ & ~new_n1738_) | ~new_n1316_ | new_n1322_)))));
  assign new_n1731_ = (((((new_n1308_ | ((new_n1632_ | ~new_n1316_ | ~new_n1322_) & ((~new_n1631_ & new_n1632_) | ~new_n1316_ | new_n1322_ | (new_n1631_ & ~new_n1632_)))) & (new_n1632_ | ~new_n1316_ | ~new_n1322_ | new_n1631_ | new_n1322_)) | ((new_n1715_ | ~new_n1316_ | ~new_n1322_) & (~new_n1316_ | new_n1322_ | (~new_n1715_ & new_n1631_ & ~new_n1632_) | (new_n1715_ & (~new_n1631_ | new_n1632_))))) & (~new_n1316_ | new_n1322_ | (new_n1631_ & ~new_n1632_) | new_n1715_ | ~new_n1322_)) | ((new_n1721_ | ~new_n1316_ | ~new_n1322_) & (~new_n1316_ | new_n1322_ | (~new_n1721_ & ~new_n1715_ & new_n1631_ & ~new_n1632_) | (new_n1721_ & (new_n1715_ | ~new_n1631_ | new_n1632_))))) & (~new_n1316_ | new_n1322_ | (~new_n1715_ & new_n1631_ & ~new_n1632_) | new_n1721_ | ~new_n1322_);
  assign new_n1732_ = ~new_n1721_ & ~new_n1715_ & new_n1631_ & ~new_n1632_;
  assign new_n1733_ = new_n1734_ & new_n1737_ & ((~P2_INSTQUEUE_REG_3__6__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_11__6__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1734_ = new_n1736_ & new_n1735_ & ((~P2_INSTQUEUE_REG_0__6__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_8__6__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1735_ = ((~P2_INSTQUEUE_REG_1__6__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_9__6__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN)) & ((~P2_INSTQUEUE_REG_2__6__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_10__6__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1736_ = ((~P2_INSTQUEUE_REG_6__6__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_14__6__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_5__6__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_13__6__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1737_ = ((~P2_INSTQUEUE_REG_7__6__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_15__6__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_4__6__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_12__6__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1738_ = new_n1739_ & new_n1742_ & ((~P2_INSTQUEUE_REG_3__5__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_11__5__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1739_ = new_n1741_ & new_n1740_ & ((~P2_INSTQUEUE_REG_0__5__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_8__5__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1740_ = ((~P2_INSTQUEUE_REG_1__5__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_9__5__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN)) & ((~P2_INSTQUEUE_REG_2__5__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_10__5__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1741_ = ((~P2_INSTQUEUE_REG_6__5__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_14__5__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_5__5__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_13__5__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1742_ = ((~P2_INSTQUEUE_REG_7__5__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_15__5__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_4__5__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_12__5__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1743_ = ~new_n1746_ ^ (new_n1744_ & ~new_n1745_);
  assign new_n1744_ = ~new_n1727_ & ~new_n1714_ & ~new_n1629_ & ~new_n1628_ & ~new_n1627_ & ~new_n1626_ & new_n1529_ & ~new_n1625_;
  assign new_n1745_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_28__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_28__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_28__SCAN_IN);
  assign new_n1746_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_29__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_29__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_29__SCAN_IN);
  assign new_n1747_ = new_n1744_ ^ ~new_n1745_;
  assign new_n1748_ = (~new_n1738_ & new_n1316_ & new_n1322_) ? (new_n1732_ | ~new_n1316_ | new_n1322_) : ((new_n1732_ | ~new_n1738_) & new_n1316_ & ~new_n1322_ & (~new_n1732_ | new_n1738_));
  assign new_n1749_ = (new_n1720_ | (new_n1726_ ^ ~new_n1727_)) & (new_n1747_ | (~new_n1731_ ^ new_n1748_));
  assign new_n1750_ = (new_n1316_ & ~new_n1322_ & (new_n1733_ | ~new_n1732_ | new_n1738_)) ^ (~new_n1751_ ^ (((~new_n1733_ & new_n1316_ & new_n1322_ & (~new_n1732_ | new_n1738_) & ~new_n1322_) | (((~new_n1733_ & new_n1316_ & new_n1322_) | (new_n1316_ & ~new_n1322_ & (new_n1733_ | ~new_n1732_ | new_n1738_) & (~new_n1733_ | (new_n1732_ & ~new_n1738_)))) & ((~new_n1738_ & new_n1316_ & new_n1322_ & ~new_n1732_ & ~new_n1322_) | (~new_n1731_ & ((~new_n1738_ & new_n1316_ & new_n1322_) | ((new_n1732_ | ~new_n1738_) & (~new_n1732_ | new_n1738_) & new_n1316_ & ~new_n1322_)))))) ^ (new_n1753_ ? (~new_n1316_ | new_n1322_) : (~new_n1316_ | ~new_n1322_))));
  assign new_n1751_ = ~new_n1752_ ^ (~new_n1746_ & new_n1744_ & ~new_n1745_);
  assign new_n1752_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_30__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_30__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_30__SCAN_IN);
  assign new_n1753_ = new_n1754_ & new_n1757_ & ((~P2_INSTQUEUE_REG_3__7__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_11__7__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1754_ = new_n1756_ & new_n1755_ & ((~P2_INSTQUEUE_REG_0__7__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_8__7__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1755_ = ((~P2_INSTQUEUE_REG_1__7__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_9__7__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN)) & ((~P2_INSTQUEUE_REG_2__7__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_10__7__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n1756_ = ((~P2_INSTQUEUE_REG_6__7__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_14__7__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_5__7__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_13__7__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1757_ = ((~P2_INSTQUEUE_REG_7__7__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUE_REG_15__7__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & ((~P2_INSTQUEUE_REG_4__7__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (~P2_INSTQUEUE_REG_12__7__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n1758_ = new_n1759_ & new_n1784_;
  assign new_n1759_ = new_n1791_ & ((new_n1760_ & new_n1364_) | new_n1785_ | (new_n1783_ & ~new_n1762_ & (new_n1768_ | ~new_n1781_)));
  assign new_n1760_ = new_n1761_ & new_n1359_;
  assign new_n1761_ = new_n1358_ & new_n1330_ & ~new_n1317_;
  assign new_n1762_ = (new_n1763_ | (P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN & (new_n1322_ | new_n1370_))) & P2_STATE2_REG_0__SCAN_IN & (new_n1322_ | new_n1370_) & (new_n1370_ | ~P2_STATE2_REG_0__SCAN_IN | (~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) | (~new_n1767_ & (~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)));
  assign new_n1763_ = ((~new_n1764_ & new_n1765_) | (~new_n1764_ & new_n1766_)) & (new_n1764_ ? ~new_n1569_ : (P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN));
  assign new_n1764_ = (~new_n1325_ | ~new_n1326_ | ~new_n1323_ | ~new_n1324_) & (~new_n1341_ | ~new_n1342_ | ~new_n1343_ | ~new_n1344_);
  assign new_n1765_ = P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n1766_ = (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & ((P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) | ((P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & ((P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))));
  assign new_n1767_ = (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) & ((P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) | ((P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & ((P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) | ((P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & ((P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))))));
  assign new_n1768_ = ~new_n1769_ & (new_n1780_ | (new_n1778_ & (new_n1771_ | ~new_n1777_ | (new_n1776_ & (~new_n1773_ | ~new_n1368_)))));
  assign new_n1769_ = ~new_n1770_ & (new_n1764_ | ~P2_STATE2_REG_0__SCAN_IN | (((~new_n1764_ & new_n1766_) | (~new_n1764_ & new_n1765_) | ((new_n1764_ | ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) & (new_n1764_ ? ~new_n1569_ : (P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)))) & ((~new_n1764_ & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) | ((new_n1764_ | ~new_n1766_) & (new_n1764_ | ~new_n1765_)) | (new_n1764_ ? new_n1569_ : (~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)))));
  assign new_n1770_ = (P2_STATE2_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN) & ((new_n1767_ & (~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ^ ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)) | (~new_n1767_ & (~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)) | ~P2_STATE2_REG_0__SCAN_IN | (new_n1343_ & new_n1344_ & new_n1341_ & new_n1342_));
  assign new_n1771_ = (((new_n1322_ | new_n1370_) & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | ((~new_n1322_ & ~new_n1370_) ? new_n1580_ : (~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) | ~new_n1370_ | ~P2_STATE2_REG_0__SCAN_IN | ((new_n1322_ | new_n1370_ | ~P2_STATE2_REG_0__SCAN_IN) & (new_n1370_ | ~P2_STATE2_REG_0__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ^ ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & (P2_STATE2_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~new_n1322_ | ~P2_STATE2_REG_0__SCAN_IN))) & (~P2_STATE2_REG_0__SCAN_IN | ((new_n1322_ | new_n1370_) & (~new_n1772_ | (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & (new_n1772_ | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) | ((new_n1370_ | (new_n1772_ & (~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) | (~new_n1772_ & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & P2_STATE2_REG_0__SCAN_IN & (new_n1322_ | ~new_n1370_))) & (new_n1322_ | new_n1370_ | ~P2_STATE2_REG_0__SCAN_IN | ((new_n1370_ | ~P2_STATE2_REG_0__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ^ ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & (P2_STATE2_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~new_n1322_ | ~P2_STATE2_REG_0__SCAN_IN)));
  assign new_n1772_ = P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n1773_ = new_n1764_ ? ~new_n1596_ : ~new_n1774_;
  assign new_n1774_ = (P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) ^ ((~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (~new_n1775_ & (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)));
  assign new_n1775_ = P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n1776_ = (~new_n1774_ | new_n1370_ | ~P2_STATE2_REG_0__SCAN_IN) & (~new_n1322_ | ~P2_STATE2_REG_0__SCAN_IN) & (P2_STATE2_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n1777_ = (P2_STATE2_REG_0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & ((P2_STATE2_REG_0__SCAN_IN & ((~new_n1322_ & ~new_n1370_) | ((~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)) | (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)))) | (~new_n1370_ & ((P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)) & (~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN))) | ~P2_STATE2_REG_0__SCAN_IN | (~new_n1322_ & new_n1370_));
  assign new_n1778_ = (new_n1322_ | new_n1370_ | new_n1779_ | ~P2_STATE2_REG_0__SCAN_IN) & (~new_n1370_ | ~P2_STATE2_REG_0__SCAN_IN | (new_n1774_ & (new_n1322_ | new_n1370_)) | (new_n1596_ & ~new_n1322_ & ~new_n1370_) | ((~new_n1774_ | new_n1370_ | ~P2_STATE2_REG_0__SCAN_IN) & (P2_STATE2_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~new_n1322_ | ~P2_STATE2_REG_0__SCAN_IN)));
  assign new_n1779_ = (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) ^ ((P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & ((P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) | ((P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & ((P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)))));
  assign new_n1780_ = (~P2_STATE2_REG_0__SCAN_IN | (~new_n1779_ & (new_n1322_ | new_n1370_))) & (P2_STATE2_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (new_n1779_ | new_n1370_ | ~P2_STATE2_REG_0__SCAN_IN);
  assign new_n1781_ = (((new_n1763_ | ((new_n1322_ | new_n1370_) & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)) & P2_STATE2_REG_0__SCAN_IN & (new_n1322_ | new_n1370_)) | new_n1370_ | ~P2_STATE2_REG_0__SCAN_IN | (~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) | (~new_n1767_ & (~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN))) & ((~P2_STATE2_REG_0__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (~new_n1370_ & P2_STATE2_REG_0__SCAN_IN & (~new_n1767_ | (P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ^ ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)) & (new_n1767_ | (P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) | (~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN))) | new_n1782_ | ~P2_STATE2_REG_0__SCAN_IN | (~new_n1322_ & ~new_n1370_));
  assign new_n1782_ = ((~new_n1764_ & new_n1765_) | (~new_n1764_ & new_n1766_) | ((new_n1764_ ? ~new_n1569_ : (P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)) & (new_n1764_ | ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN))) & (((new_n1764_ | ~new_n1765_) & (new_n1764_ | ~new_n1766_)) | (new_n1764_ ? new_n1569_ : (~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)) | (~new_n1764_ & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN));
  assign new_n1783_ = new_n1364_ & new_n1367_ & new_n1784_ & ~new_n1345_ & ~new_n1335_ & ~new_n1350_;
  assign new_n1784_ = ~new_n1330_ & new_n1317_;
  assign new_n1785_ = new_n1788_ & ~new_n1790_ & ((new_n1786_ & new_n1322_) | (new_n1787_ & ~new_n1322_ & ~new_n1370_));
  assign new_n1786_ = ~new_n1335_ & ~new_n1317_ & ~new_n1330_ & new_n1350_ & new_n1370_ & new_n1345_ & ~new_n1367_;
  assign new_n1787_ = new_n1330_ & new_n1377_ & new_n1350_ & new_n1356_;
  assign new_n1788_ = ((~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) | (~new_n1767_ & (~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN))) & (~new_n1789_ | ~new_n1779_ | (new_n1767_ ^ (~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ^ ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)));
  assign new_n1789_ = ((P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) ^ ((~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | ((~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)))) & ((P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) ^ (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN));
  assign new_n1790_ = READY12_REG_SCAN_IN & READY21_REG_SCAN_IN;
  assign new_n1791_ = new_n1792_ & P2_STATE2_REG_0__SCAN_IN;
  assign new_n1792_ = P2_STATE2_REG_2__SCAN_IN & ~P2_STATE2_REG_1__SCAN_IN;
  assign new_n1793_ = ~new_n1794_ & new_n4475_ & new_n4491_ & ~new_n2041_ & ~new_n4506_ & new_n2499_ & new_n4468_;
  assign new_n1794_ = new_n1957_ & ((new_n2030_ & (~new_n2038_ | ((new_n2039_ | (~new_n1795_ & P2_INSTADDRPOINTER_REG_25__SCAN_IN)) & new_n2034_ & (~new_n1795_ | P2_INSTADDRPOINTER_REG_25__SCAN_IN)))) | ~new_n2040_ | (~new_n2030_ & new_n2038_ & ((~new_n2039_ & (new_n1795_ | ~P2_INSTADDRPOINTER_REG_25__SCAN_IN)) | ~new_n2034_ | (new_n1795_ & ~P2_INSTADDRPOINTER_REG_25__SCAN_IN))));
  assign new_n1795_ = new_n1950_ & ((new_n1955_ & (~new_n1952_ | (new_n1951_ & (new_n1796_ | ~new_n1937_)))) | new_n1945_ | new_n1956_);
  assign new_n1796_ = new_n1928_ & (new_n1921_ | (new_n1936_ & (~new_n1933_ | new_n1930_ | (~new_n1932_ & (new_n1797_ | new_n1927_)))));
  assign new_n1797_ = new_n1919_ & (~new_n1912_ | (new_n1911_ & (~new_n1904_ | (~new_n1798_ & (new_n1880_ | (~new_n1881_ & ~new_n1884_))))));
  assign new_n1798_ = P2_INSTADDRPOINTER_REG_7__SCAN_IN & ((new_n1799_ & new_n1534_) | ((new_n1870_ | new_n1878_) & ~new_n1534_ & (~new_n1870_ | ~new_n1878_)));
  assign new_n1799_ = ~new_n1800_ ^ (~new_n1865_ & ~new_n1860_ & ~new_n1855_ & new_n1820_ & new_n1849_);
  assign new_n1800_ = new_n1322_ ? new_n1534_ : (new_n1812_ & new_n1815_ & new_n1801_ & new_n1807_);
  assign new_n1801_ = (~new_n1802_ | ~P2_INSTQUEUE_REG_10__7__SCAN_IN) & (~new_n1804_ | ~P2_INSTQUEUE_REG_1__7__SCAN_IN) & (~new_n1805_ | ~P2_INSTQUEUE_REG_7__7__SCAN_IN) & (~new_n1806_ | ~P2_INSTQUEUE_REG_13__7__SCAN_IN);
  assign new_n1802_ = new_n1413_ & ~new_n1803_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_)) & (new_n1387_ ^ (~new_n1383_ & ~new_n1386_));
  assign new_n1803_ = (~new_n1390_ & (~new_n1328_ | ~new_n1388_)) ^ (new_n1391_ | ~new_n1392_);
  assign new_n1804_ = ~new_n1413_ & new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ ^ (~new_n1383_ & ~new_n1386_));
  assign new_n1805_ = new_n1413_ & new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1806_ = ~new_n1413_ & new_n1803_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_)) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1807_ = (~new_n1809_ | ~P2_INSTQUEUE_REG_0__7__SCAN_IN) & (~new_n1808_ | ~P2_INSTQUEUE_REG_3__7__SCAN_IN) & (~new_n1811_ | ~P2_INSTQUEUE_REG_5__7__SCAN_IN) & (~new_n1810_ | ~P2_INSTQUEUE_REG_11__7__SCAN_IN);
  assign new_n1808_ = new_n1413_ & new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ ^ (~new_n1383_ & ~new_n1386_));
  assign new_n1809_ = ~new_n1413_ & ~new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ ^ (~new_n1383_ & ~new_n1386_));
  assign new_n1810_ = new_n1413_ & new_n1803_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_)) & (new_n1387_ ^ (~new_n1383_ & ~new_n1386_));
  assign new_n1811_ = ~new_n1413_ & new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1812_ = (~P2_INSTQUEUE_REG_6__7__SCAN_IN | new_n1813_ | ~new_n1814_ | ~new_n1413_ | new_n1803_) & (~P2_INSTQUEUE_REG_8__7__SCAN_IN | new_n1413_ | new_n1803_ | ~new_n1813_ | new_n1814_) & (~P2_INSTQUEUE_REG_14__7__SCAN_IN | ~new_n1813_ | ~new_n1814_ | ~new_n1413_ | new_n1803_) & (~P2_INSTQUEUE_REG_4__7__SCAN_IN | new_n1413_ | new_n1803_ | new_n1813_ | ~new_n1814_);
  assign new_n1813_ = new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_));
  assign new_n1814_ = new_n1387_ ^ ~new_n1410_;
  assign new_n1815_ = (~new_n1817_ | ~P2_INSTQUEUE_REG_15__7__SCAN_IN) & (~new_n1816_ | ~P2_INSTQUEUE_REG_2__7__SCAN_IN) & (~new_n1819_ | ~P2_INSTQUEUE_REG_9__7__SCAN_IN) & (~new_n1818_ | ~P2_INSTQUEUE_REG_12__7__SCAN_IN);
  assign new_n1816_ = new_n1413_ & ~new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ ^ (~new_n1383_ & ~new_n1386_));
  assign new_n1817_ = new_n1413_ & new_n1803_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_)) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1818_ = ~new_n1413_ & ~new_n1803_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_)) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1819_ = ~new_n1413_ & new_n1803_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_)) & (new_n1387_ ^ (~new_n1383_ & ~new_n1386_));
  assign new_n1820_ = (~new_n1837_ | ~new_n1841_ | ~new_n1842_) & ((new_n1322_ & ~new_n1596_) | new_n1848_ | (~new_n1322_ & (~new_n1821_ | ~new_n1828_)));
  assign new_n1821_ = ~new_n1823_ & ~new_n1824_ & ~new_n1822_ & (~new_n1809_ | ~P2_INSTQUEUE_REG_0__1__SCAN_IN) & new_n1825_ & ~new_n1826_ & ~new_n1827_;
  assign new_n1822_ = P2_INSTQUEUE_REG_1__1__SCAN_IN & ~new_n1413_ & new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ ^ (~new_n1383_ & ~new_n1386_));
  assign new_n1823_ = P2_INSTQUEUE_REG_5__1__SCAN_IN & ~new_n1413_ & new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1824_ = P2_INSTQUEUE_REG_11__1__SCAN_IN & new_n1413_ & new_n1803_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_)) & (new_n1387_ ^ (~new_n1383_ & ~new_n1386_));
  assign new_n1825_ = (~P2_INSTQUEUE_REG_8__1__SCAN_IN | new_n1413_ | new_n1803_ | (new_n1327_ & (new_n1383_ | (~new_n1386_ & ~new_n1387_))) | (~new_n1327_ & ~new_n1383_ & (new_n1386_ | new_n1387_)) | (~new_n1387_ ^ (~new_n1383_ & ~new_n1386_))) & (~P2_INSTQUEUE_REG_9__1__SCAN_IN | new_n1413_ | ~new_n1803_ | (new_n1327_ & (new_n1383_ | (~new_n1386_ & ~new_n1387_))) | (~new_n1327_ & ~new_n1383_ & (new_n1386_ | new_n1387_)) | (~new_n1387_ ^ (~new_n1383_ & ~new_n1386_)));
  assign new_n1826_ = P2_INSTQUEUE_REG_6__1__SCAN_IN & new_n1413_ & ~new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1827_ = P2_INSTQUEUE_REG_7__1__SCAN_IN & new_n1413_ & new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1828_ = ~new_n1831_ & ~new_n1832_ & ~new_n1829_ & ~new_n1830_ & ~new_n1833_ & ~new_n1834_ & ~new_n1835_ & ~new_n1836_;
  assign new_n1829_ = P2_INSTQUEUE_REG_2__1__SCAN_IN & new_n1413_ & ~new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ ^ (~new_n1383_ & ~new_n1386_));
  assign new_n1830_ = P2_INSTQUEUE_REG_13__1__SCAN_IN & ~new_n1413_ & new_n1803_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_)) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1831_ = P2_INSTQUEUE_REG_10__1__SCAN_IN & new_n1413_ & ~new_n1803_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_)) & (new_n1387_ ^ (~new_n1383_ & ~new_n1386_));
  assign new_n1832_ = P2_INSTQUEUE_REG_12__1__SCAN_IN & ~new_n1413_ & ~new_n1803_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_)) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1833_ = P2_INSTQUEUE_REG_4__1__SCAN_IN & ~new_n1413_ & ~new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1834_ = P2_INSTQUEUE_REG_3__1__SCAN_IN & new_n1413_ & new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ ^ (~new_n1383_ & ~new_n1386_));
  assign new_n1835_ = P2_INSTQUEUE_REG_14__1__SCAN_IN & new_n1413_ & ~new_n1803_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_)) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1836_ = P2_INSTQUEUE_REG_15__1__SCAN_IN & new_n1413_ & new_n1803_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_)) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1837_ = new_n1839_ & (~new_n1802_ | ~P2_INSTQUEUE_REG_10__2__SCAN_IN) & (~new_n1817_ | ~P2_INSTQUEUE_REG_15__2__SCAN_IN) & ~new_n1840_ & (~new_n1838_ | ~P2_INSTQUEUE_REG_14__2__SCAN_IN);
  assign new_n1838_ = new_n1413_ & ~new_n1803_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_)) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1839_ = ~new_n1322_ & (~P2_INSTQUEUE_REG_2__2__SCAN_IN | ~new_n1413_ | new_n1803_ | (new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) | (~new_n1387_ ^ (~new_n1383_ & ~new_n1386_)));
  assign new_n1840_ = P2_INSTQUEUE_REG_9__2__SCAN_IN & ~new_n1413_ & new_n1803_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_)) & (new_n1387_ ^ (~new_n1383_ & ~new_n1386_));
  assign new_n1841_ = (~new_n1818_ | ~P2_INSTQUEUE_REG_12__2__SCAN_IN) & (~new_n1806_ | ~P2_INSTQUEUE_REG_13__2__SCAN_IN) & (~new_n1809_ | ~P2_INSTQUEUE_REG_0__2__SCAN_IN);
  assign new_n1842_ = new_n1844_ & new_n1845_ & ~new_n1846_ & ~new_n1847_ & (~new_n1843_ | ~P2_INSTQUEUE_REG_4__2__SCAN_IN) & (~new_n1811_ | ~P2_INSTQUEUE_REG_5__2__SCAN_IN);
  assign new_n1843_ = ~new_n1413_ & ~new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1844_ = (~P2_INSTQUEUE_REG_8__2__SCAN_IN | new_n1413_ | new_n1803_ | (new_n1327_ & (new_n1383_ | (~new_n1386_ & ~new_n1387_))) | (~new_n1327_ & ~new_n1383_ & (new_n1386_ | new_n1387_)) | (~new_n1387_ ^ (~new_n1383_ & ~new_n1386_))) & (~P2_INSTQUEUE_REG_7__2__SCAN_IN | ~new_n1413_ | ~new_n1803_ | (new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) | (~new_n1387_ & ~new_n1383_ & ~new_n1386_) | (new_n1387_ & (new_n1383_ | new_n1386_)));
  assign new_n1845_ = (~P2_INSTQUEUE_REG_11__2__SCAN_IN | ~new_n1413_ | ~new_n1803_ | (new_n1327_ & (new_n1383_ | (~new_n1386_ & ~new_n1387_))) | (~new_n1327_ & ~new_n1383_ & (new_n1386_ | new_n1387_)) | (~new_n1387_ ^ (~new_n1383_ & ~new_n1386_))) & (~P2_INSTQUEUE_REG_3__2__SCAN_IN | ~new_n1413_ | ~new_n1803_ | (new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) | (~new_n1387_ ^ (~new_n1383_ & ~new_n1386_)));
  assign new_n1846_ = P2_INSTQUEUE_REG_1__2__SCAN_IN & ~new_n1413_ & new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ ^ (~new_n1383_ & ~new_n1386_));
  assign new_n1847_ = P2_INSTQUEUE_REG_6__2__SCAN_IN & new_n1413_ & ~new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1848_ = ~new_n1580_ & new_n1322_ & ~new_n1587_;
  assign new_n1849_ = (~new_n1322_ | ~new_n1607_) & (~new_n1851_ | ~new_n1852_ | ~new_n1853_ | ~new_n1850_ | new_n1322_ | (new_n1818_ & P2_INSTQUEUE_REG_12__3__SCAN_IN));
  assign new_n1850_ = (~new_n1810_ | ~P2_INSTQUEUE_REG_11__3__SCAN_IN) & (~new_n1808_ | ~P2_INSTQUEUE_REG_3__3__SCAN_IN) & (~new_n1838_ | ~P2_INSTQUEUE_REG_14__3__SCAN_IN) & (~new_n1805_ | ~P2_INSTQUEUE_REG_7__3__SCAN_IN);
  assign new_n1851_ = (~new_n1817_ | ~P2_INSTQUEUE_REG_15__3__SCAN_IN) & (~new_n1806_ | ~P2_INSTQUEUE_REG_13__3__SCAN_IN) & (~new_n1819_ | ~P2_INSTQUEUE_REG_9__3__SCAN_IN);
  assign new_n1852_ = (~P2_INSTQUEUE_REG_10__3__SCAN_IN | ~new_n1813_ | new_n1814_ | ~new_n1413_ | new_n1803_) & (~P2_INSTQUEUE_REG_1__3__SCAN_IN | new_n1813_ | new_n1814_ | new_n1413_ | ~new_n1803_) & (~P2_INSTQUEUE_REG_8__3__SCAN_IN | new_n1413_ | new_n1803_ | ~new_n1813_ | new_n1814_) & (~P2_INSTQUEUE_REG_2__3__SCAN_IN | new_n1813_ | new_n1814_ | ~new_n1413_ | new_n1803_);
  assign new_n1853_ = (~new_n1811_ | ~P2_INSTQUEUE_REG_5__3__SCAN_IN) & (~new_n1843_ | ~P2_INSTQUEUE_REG_4__3__SCAN_IN) & (~new_n1809_ | ~P2_INSTQUEUE_REG_0__3__SCAN_IN) & (~new_n1854_ | ~P2_INSTQUEUE_REG_6__3__SCAN_IN);
  assign new_n1854_ = new_n1413_ & ~new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_));
  assign new_n1855_ = new_n1322_ ? new_n1569_ : (new_n1858_ & new_n1859_ & new_n1856_ & new_n1857_);
  assign new_n1856_ = (~new_n1802_ | ~P2_INSTQUEUE_REG_10__4__SCAN_IN) & (~new_n1804_ | ~P2_INSTQUEUE_REG_1__4__SCAN_IN) & (~new_n1805_ | ~P2_INSTQUEUE_REG_7__4__SCAN_IN) & (~new_n1806_ | ~P2_INSTQUEUE_REG_13__4__SCAN_IN);
  assign new_n1857_ = (~new_n1809_ | ~P2_INSTQUEUE_REG_0__4__SCAN_IN) & (~new_n1808_ | ~P2_INSTQUEUE_REG_3__4__SCAN_IN) & (~new_n1811_ | ~P2_INSTQUEUE_REG_5__4__SCAN_IN) & (~new_n1810_ | ~P2_INSTQUEUE_REG_11__4__SCAN_IN);
  assign new_n1858_ = (~P2_INSTQUEUE_REG_6__4__SCAN_IN | new_n1813_ | ~new_n1814_ | ~new_n1413_ | new_n1803_) & (~P2_INSTQUEUE_REG_8__4__SCAN_IN | new_n1413_ | new_n1803_ | ~new_n1813_ | new_n1814_) & (~P2_INSTQUEUE_REG_14__4__SCAN_IN | ~new_n1813_ | ~new_n1814_ | ~new_n1413_ | new_n1803_) & (~P2_INSTQUEUE_REG_4__4__SCAN_IN | new_n1413_ | new_n1803_ | new_n1813_ | ~new_n1814_);
  assign new_n1859_ = (~new_n1817_ | ~P2_INSTQUEUE_REG_15__4__SCAN_IN) & (~new_n1816_ | ~P2_INSTQUEUE_REG_2__4__SCAN_IN) & (~new_n1819_ | ~P2_INSTQUEUE_REG_9__4__SCAN_IN) & (~new_n1818_ | ~P2_INSTQUEUE_REG_12__4__SCAN_IN);
  assign new_n1860_ = new_n1322_ ? new_n1560_ : (new_n1863_ & new_n1864_ & new_n1861_ & new_n1862_);
  assign new_n1861_ = (~new_n1802_ | ~P2_INSTQUEUE_REG_10__5__SCAN_IN) & (~new_n1804_ | ~P2_INSTQUEUE_REG_1__5__SCAN_IN) & (~new_n1805_ | ~P2_INSTQUEUE_REG_7__5__SCAN_IN) & (~new_n1806_ | ~P2_INSTQUEUE_REG_13__5__SCAN_IN);
  assign new_n1862_ = (~new_n1809_ | ~P2_INSTQUEUE_REG_0__5__SCAN_IN) & (~new_n1808_ | ~P2_INSTQUEUE_REG_3__5__SCAN_IN) & (~new_n1811_ | ~P2_INSTQUEUE_REG_5__5__SCAN_IN) & (~new_n1810_ | ~P2_INSTQUEUE_REG_11__5__SCAN_IN);
  assign new_n1863_ = (~P2_INSTQUEUE_REG_6__5__SCAN_IN | new_n1813_ | ~new_n1814_ | ~new_n1413_ | new_n1803_) & (~P2_INSTQUEUE_REG_8__5__SCAN_IN | new_n1413_ | new_n1803_ | ~new_n1813_ | new_n1814_) & (~P2_INSTQUEUE_REG_14__5__SCAN_IN | ~new_n1813_ | ~new_n1814_ | ~new_n1413_ | new_n1803_) & (~P2_INSTQUEUE_REG_4__5__SCAN_IN | new_n1413_ | new_n1803_ | new_n1813_ | ~new_n1814_);
  assign new_n1864_ = (~new_n1817_ | ~P2_INSTQUEUE_REG_15__5__SCAN_IN) & (~new_n1816_ | ~P2_INSTQUEUE_REG_2__5__SCAN_IN) & (~new_n1819_ | ~P2_INSTQUEUE_REG_9__5__SCAN_IN) & (~new_n1818_ | ~P2_INSTQUEUE_REG_12__5__SCAN_IN);
  assign new_n1865_ = new_n1322_ ? new_n1551_ : (new_n1868_ & new_n1869_ & new_n1866_ & new_n1867_);
  assign new_n1866_ = (~new_n1802_ | ~P2_INSTQUEUE_REG_10__6__SCAN_IN) & (~new_n1804_ | ~P2_INSTQUEUE_REG_1__6__SCAN_IN) & (~new_n1805_ | ~P2_INSTQUEUE_REG_7__6__SCAN_IN) & (~new_n1806_ | ~P2_INSTQUEUE_REG_13__6__SCAN_IN);
  assign new_n1867_ = (~new_n1809_ | ~P2_INSTQUEUE_REG_0__6__SCAN_IN) & (~new_n1808_ | ~P2_INSTQUEUE_REG_3__6__SCAN_IN) & (~new_n1811_ | ~P2_INSTQUEUE_REG_5__6__SCAN_IN) & (~new_n1810_ | ~P2_INSTQUEUE_REG_11__6__SCAN_IN);
  assign new_n1868_ = (~P2_INSTQUEUE_REG_6__6__SCAN_IN | new_n1813_ | ~new_n1814_ | ~new_n1413_ | new_n1803_) & (~P2_INSTQUEUE_REG_8__6__SCAN_IN | new_n1413_ | new_n1803_ | ~new_n1813_ | new_n1814_) & (~P2_INSTQUEUE_REG_14__6__SCAN_IN | ~new_n1813_ | ~new_n1814_ | ~new_n1413_ | new_n1803_) & (~P2_INSTQUEUE_REG_4__6__SCAN_IN | new_n1413_ | new_n1803_ | new_n1813_ | ~new_n1814_);
  assign new_n1869_ = (~new_n1817_ | ~P2_INSTQUEUE_REG_15__6__SCAN_IN) & (~new_n1816_ | ~P2_INSTQUEUE_REG_2__6__SCAN_IN) & (~new_n1819_ | ~P2_INSTQUEUE_REG_9__6__SCAN_IN) & (~new_n1818_ | ~P2_INSTQUEUE_REG_12__6__SCAN_IN);
  assign new_n1870_ = new_n1871_ & ~new_n1876_;
  assign new_n1871_ = ~new_n1874_ & new_n1872_ & ~new_n1873_ & (new_n1330_ ? ~P2_EBX_REG_4__SCAN_IN : new_n1782_) & (~new_n1330_ | ~P2_EBX_REG_5__SCAN_IN) & (new_n1875_ | new_n1330_);
  assign new_n1872_ = (~new_n1330_ | (~P2_EBX_REG_0__SCAN_IN & ~P2_EBX_REG_1__SCAN_IN)) & (((~new_n1587_ | ~new_n1764_) & (new_n1764_ | new_n1772_) & (new_n1764_ | ~new_n1775_)) | new_n1330_ | (new_n1775_ & ~new_n1764_ & ~new_n1772_));
  assign new_n1873_ = new_n1330_ ? P2_EBX_REG_2__SCAN_IN : (new_n1764_ ? new_n1596_ : new_n1774_);
  assign new_n1874_ = new_n1330_ ? P2_EBX_REG_3__SCAN_IN : (new_n1764_ ? new_n1607_ : ~new_n1779_);
  assign new_n1875_ = (new_n1560_ & new_n1764_) ? (((~new_n1764_ & new_n1766_) | (~new_n1764_ & new_n1765_)) & (new_n1764_ ? ~new_n1569_ : (P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN))) : ((new_n1764_ | ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) & (((new_n1764_ | ~new_n1766_) & (new_n1764_ | ~new_n1765_)) | (new_n1764_ ? new_n1569_ : (~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN))));
  assign new_n1876_ = (~new_n1330_ | P2_EBX_REG_6__SCAN_IN) & ((new_n1551_ & new_n1764_ & (new_n1877_ | (new_n1560_ & new_n1764_))) | new_n1330_ | ((~new_n1551_ | ~new_n1764_) & ~new_n1877_ & (~new_n1560_ | ~new_n1764_)));
  assign new_n1877_ = (((new_n1764_ | ~new_n1765_) & (new_n1764_ | ~new_n1766_)) | (new_n1764_ ? new_n1569_ : (~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN))) & (new_n1764_ | ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  assign new_n1878_ = (new_n1879_ | new_n1330_ | ~new_n1534_ | ~new_n1764_) & (~new_n1330_ | ~P2_EBX_REG_7__SCAN_IN) & (~new_n1879_ | new_n1330_ | (new_n1534_ & new_n1764_));
  assign new_n1879_ = (~new_n1551_ | ~new_n1764_) & (~new_n1560_ | ~new_n1764_) & ((~new_n1764_ & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) | (((~new_n1764_ & new_n1765_) | (~new_n1764_ & new_n1766_)) & (new_n1764_ ? ~new_n1569_ : (P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN))));
  assign new_n1880_ = ~P2_INSTADDRPOINTER_REG_7__SCAN_IN & (~new_n1799_ | ~new_n1534_) & ((~new_n1870_ & ~new_n1878_) | new_n1534_ | (new_n1870_ & new_n1878_));
  assign new_n1881_ = P2_INSTADDRPOINTER_REG_6__SCAN_IN & (new_n1534_ ? (new_n1882_ ^ ~new_n1865_) : new_n1883_);
  assign new_n1882_ = ~new_n1860_ & ~new_n1855_ & new_n1820_ & new_n1849_;
  assign new_n1883_ = new_n1871_ ^ ~new_n1876_;
  assign new_n1884_ = ~new_n1885_ & ((~new_n1886_ & P2_INSTADDRPOINTER_REG_5__SCAN_IN) | ((~new_n1886_ | P2_INSTADDRPOINTER_REG_5__SCAN_IN) & ((~new_n1890_ & P2_INSTADDRPOINTER_REG_4__SCAN_IN) | ((~new_n1903_ | (~new_n1892_ & P2_INSTADDRPOINTER_REG_3__SCAN_IN)) & (~new_n1890_ | P2_INSTADDRPOINTER_REG_4__SCAN_IN) & (~new_n1892_ | P2_INSTADDRPOINTER_REG_3__SCAN_IN)))));
  assign new_n1885_ = ~P2_INSTADDRPOINTER_REG_6__SCAN_IN & (~new_n1883_ | new_n1534_) & (~new_n1534_ | (~new_n1865_ & ~new_n1860_ & ~new_n1855_ & new_n1820_ & new_n1849_) | (new_n1865_ & (new_n1860_ | new_n1855_ | ~new_n1820_ | ~new_n1849_)));
  assign new_n1886_ = ~new_n1887_ & (~new_n1534_ | (~new_n1860_ & ~new_n1855_ & new_n1820_ & new_n1849_) | (new_n1860_ & (new_n1855_ | ~new_n1820_ | ~new_n1849_)));
  assign new_n1887_ = ((new_n1888_ & (new_n1330_ ? ~P2_EBX_REG_4__SCAN_IN : new_n1782_)) | (new_n1330_ ? ~P2_EBX_REG_5__SCAN_IN : new_n1875_)) & ~new_n1534_ & (~new_n1888_ | (new_n1330_ ? P2_EBX_REG_4__SCAN_IN : ~new_n1782_) | (new_n1330_ & P2_EBX_REG_5__SCAN_IN) | (~new_n1875_ & ~new_n1330_));
  assign new_n1888_ = new_n1889_ & ~new_n1874_;
  assign new_n1889_ = new_n1872_ & ~new_n1873_;
  assign new_n1890_ = new_n1534_ ? (new_n1855_ ^ (new_n1820_ & new_n1849_)) : ~new_n1891_;
  assign new_n1891_ = new_n1888_ ^ (new_n1330_ ? ~P2_EBX_REG_4__SCAN_IN : new_n1782_);
  assign new_n1892_ = (~P2_INSTADDRPOINTER_REG_2__SCAN_IN | (new_n1534_ ? ~new_n1893_ : ~new_n1902_)) & ((~new_n1900_ & (~new_n1894_ | ~P2_INSTADDRPOINTER_REG_1__SCAN_IN)) | (~new_n1894_ & ~P2_INSTADDRPOINTER_REG_1__SCAN_IN) | (~P2_INSTADDRPOINTER_REG_2__SCAN_IN & (~new_n1893_ | ~new_n1534_) & (~new_n1902_ | new_n1534_)));
  assign new_n1893_ = (~new_n1848_ & (new_n1322_ | (new_n1821_ & new_n1828_))) ^ ((new_n1322_ & ~new_n1596_) | (new_n1837_ & new_n1841_ & new_n1842_));
  assign new_n1894_ = new_n1899_ & (~new_n1534_ | (new_n1322_ & new_n1580_) | (~new_n1322_ & (~new_n1897_ | ~new_n1898_ | ~new_n1895_ | ~new_n1896_)));
  assign new_n1895_ = (~new_n1809_ | ~P2_INSTQUEUE_REG_0__0__SCAN_IN) & (~new_n1804_ | ~P2_INSTQUEUE_REG_1__0__SCAN_IN) & (~new_n1854_ | ~P2_INSTQUEUE_REG_6__0__SCAN_IN) & (~new_n1806_ | ~P2_INSTQUEUE_REG_13__0__SCAN_IN);
  assign new_n1896_ = (~P2_INSTQUEUE_REG_8__0__SCAN_IN | new_n1413_ | new_n1803_ | ~new_n1813_ | new_n1814_) & (~P2_INSTQUEUE_REG_9__0__SCAN_IN | ~new_n1813_ | new_n1814_ | new_n1413_ | ~new_n1803_) & (~P2_INSTQUEUE_REG_7__0__SCAN_IN | ~new_n1413_ | ~new_n1803_ | new_n1813_ | ~new_n1814_) & (~P2_INSTQUEUE_REG_3__0__SCAN_IN | ~new_n1413_ | ~new_n1803_ | new_n1813_ | new_n1814_);
  assign new_n1897_ = (~new_n1838_ | ~P2_INSTQUEUE_REG_14__0__SCAN_IN) & (~new_n1816_ | ~P2_INSTQUEUE_REG_2__0__SCAN_IN) & (~new_n1818_ | ~P2_INSTQUEUE_REG_12__0__SCAN_IN) & (~new_n1802_ | ~P2_INSTQUEUE_REG_10__0__SCAN_IN);
  assign new_n1898_ = (~new_n1843_ | ~P2_INSTQUEUE_REG_4__0__SCAN_IN) & (~new_n1811_ | ~P2_INSTQUEUE_REG_5__0__SCAN_IN) & (~new_n1817_ | ~P2_INSTQUEUE_REG_15__0__SCAN_IN) & (~new_n1810_ | ~P2_INSTQUEUE_REG_11__0__SCAN_IN);
  assign new_n1899_ = P2_INSTADDRPOINTER_REG_0__SCAN_IN & ((~new_n1330_ & (new_n1764_ | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (new_n1764_ ? ~new_n1580_ : (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))) | new_n1534_ | (new_n1330_ & P2_EBX_REG_0__SCAN_IN));
  assign new_n1900_ = new_n1534_ ? ((~new_n1587_ | ~new_n1322_ | ~new_n1580_) & (new_n1580_ | ~new_n1322_ | new_n1587_) & (new_n1322_ | (new_n1821_ & new_n1828_))) : new_n1901_;
  assign new_n1901_ = ~new_n1872_ & (~P2_EBX_REG_1__SCAN_IN | ~new_n1330_ | ~P2_EBX_REG_0__SCAN_IN);
  assign new_n1902_ = new_n1872_ ^ ~new_n1873_;
  assign new_n1903_ = (~new_n1534_ | (new_n1820_ & new_n1849_) | (~new_n1820_ & ~new_n1849_)) & ((~new_n1889_ & new_n1874_) | new_n1534_ | (new_n1889_ & ~new_n1874_));
  assign new_n1904_ = (new_n1906_ | P2_INSTADDRPOINTER_REG_9__SCAN_IN) & (P2_INSTADDRPOINTER_REG_8__SCAN_IN | (new_n1534_ ? new_n1905_ : new_n1910_));
  assign new_n1905_ = ~new_n1800_ & ~new_n1865_ & ~new_n1860_ & ~new_n1855_ & new_n1820_ & new_n1849_;
  assign new_n1906_ = ((~new_n1907_ & ~new_n1908_) | (~new_n1909_ & new_n1870_ & new_n1878_)) & ~new_n1534_ & (new_n1908_ | new_n1909_ | ~new_n1870_ | ~new_n1878_);
  assign new_n1907_ = new_n1879_ & ~new_n1330_ & (~new_n1534_ | ~new_n1764_);
  assign new_n1908_ = new_n1330_ & P2_EBX_REG_9__SCAN_IN;
  assign new_n1909_ = new_n1330_ & P2_EBX_REG_8__SCAN_IN;
  assign new_n1910_ = (new_n1870_ & new_n1878_) ? new_n1909_ : (~new_n1907_ & ~new_n1909_);
  assign new_n1911_ = (~new_n1906_ | ~P2_INSTADDRPOINTER_REG_9__SCAN_IN) & ((~new_n1906_ & ~P2_INSTADDRPOINTER_REG_9__SCAN_IN) | ~P2_INSTADDRPOINTER_REG_8__SCAN_IN | (~new_n1905_ & new_n1534_) | (~new_n1910_ & ~new_n1534_));
  assign new_n1912_ = (P2_INSTADDRPOINTER_REG_11__SCAN_IN | (~new_n1917_ & ~new_n1913_ & ~new_n1534_)) & (P2_INSTADDRPOINTER_REG_10__SCAN_IN | (new_n1918_ & ~new_n1534_));
  assign new_n1913_ = ~new_n1916_ & new_n1914_ & new_n1915_;
  assign new_n1914_ = ~new_n1908_ & ~new_n1909_ & new_n1870_ & new_n1878_;
  assign new_n1915_ = (~new_n1330_ | ~P2_EBX_REG_10__SCAN_IN) & (~new_n1879_ | new_n1330_ | (new_n1534_ & new_n1764_));
  assign new_n1916_ = new_n1330_ & P2_EBX_REG_11__SCAN_IN;
  assign new_n1917_ = (~new_n1914_ | ~new_n1915_) & (new_n1907_ | new_n1916_);
  assign new_n1918_ = new_n1914_ ^ new_n1915_;
  assign new_n1919_ = ((~P2_INSTADDRPOINTER_REG_11__SCAN_IN & (new_n1917_ | new_n1913_ | new_n1534_)) | ~P2_INSTADDRPOINTER_REG_10__SCAN_IN | ~new_n1918_ | new_n1534_) & (~P2_INSTADDRPOINTER_REG_12__SCAN_IN | (~new_n1913_ & ~new_n1920_) | new_n1534_ | (new_n1913_ & new_n1920_)) & (~P2_INSTADDRPOINTER_REG_11__SCAN_IN | new_n1917_ | new_n1913_ | new_n1534_);
  assign new_n1920_ = (~new_n1330_ | ~P2_EBX_REG_12__SCAN_IN) & (~new_n1879_ | new_n1330_ | (new_n1534_ & new_n1764_));
  assign new_n1921_ = ~new_n1922_ & ~P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign new_n1922_ = (new_n1923_ | new_n1926_) & ~new_n1534_ & (~new_n1923_ | ~new_n1926_);
  assign new_n1923_ = (~new_n1330_ | ~P2_EBX_REG_15__SCAN_IN) & new_n1924_ & new_n1925_ & (~new_n1330_ | ~P2_EBX_REG_13__SCAN_IN);
  assign new_n1924_ = ~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_14__SCAN_IN);
  assign new_n1925_ = new_n1920_ & ~new_n1916_ & new_n1915_ & ~new_n1908_ & ~new_n1909_ & new_n1878_ & new_n1871_ & ~new_n1876_;
  assign new_n1926_ = ~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_16__SCAN_IN);
  assign new_n1927_ = ~P2_INSTADDRPOINTER_REG_12__SCAN_IN & ((~new_n1913_ & ~new_n1920_) | new_n1534_ | (new_n1913_ & new_n1920_));
  assign new_n1928_ = (~new_n1922_ | ~P2_INSTADDRPOINTER_REG_16__SCAN_IN) & (~new_n1929_ | ~P2_INSTADDRPOINTER_REG_17__SCAN_IN);
  assign new_n1929_ = ((new_n1923_ & ~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_16__SCAN_IN)) | (~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_17__SCAN_IN))) & ~new_n1534_ & ((new_n1330_ & P2_EBX_REG_17__SCAN_IN) | ~new_n1923_ | new_n1907_ | (new_n1330_ & P2_EBX_REG_16__SCAN_IN));
  assign new_n1930_ = ~new_n1931_ & ~P2_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign new_n1931_ = ~new_n1534_ & (new_n1925_ | ~new_n1330_ | ~P2_EBX_REG_13__SCAN_IN) & ~new_n1907_ & (~new_n1925_ | (new_n1330_ & P2_EBX_REG_13__SCAN_IN));
  assign new_n1932_ = new_n1931_ & P2_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign new_n1933_ = (new_n1935_ | P2_INSTADDRPOINTER_REG_14__SCAN_IN) & (new_n1934_ | P2_INSTADDRPOINTER_REG_15__SCAN_IN);
  assign new_n1934_ = ~new_n1534_ & (~new_n1330_ | ~P2_EBX_REG_15__SCAN_IN | (new_n1924_ & new_n1925_ & (~new_n1330_ | ~P2_EBX_REG_13__SCAN_IN))) & ~new_n1907_ & ((new_n1330_ & P2_EBX_REG_15__SCAN_IN) | ~new_n1924_ | ~new_n1925_ | (new_n1330_ & P2_EBX_REG_13__SCAN_IN));
  assign new_n1935_ = (new_n1924_ | (new_n1925_ & (~new_n1330_ | ~P2_EBX_REG_13__SCAN_IN))) & ~new_n1534_ & (~new_n1924_ | ~new_n1925_ | (new_n1330_ & P2_EBX_REG_13__SCAN_IN));
  assign new_n1936_ = (~new_n1934_ | ~P2_INSTADDRPOINTER_REG_15__SCAN_IN) & ((~new_n1934_ & ~P2_INSTADDRPOINTER_REG_15__SCAN_IN) | ~new_n1935_ | ~P2_INSTADDRPOINTER_REG_14__SCAN_IN);
  assign new_n1937_ = new_n1938_ & (new_n1941_ | P2_INSTADDRPOINTER_REG_19__SCAN_IN) & (P2_INSTADDRPOINTER_REG_20__SCAN_IN | (new_n1943_ & ~new_n1534_));
  assign new_n1938_ = (new_n1929_ | P2_INSTADDRPOINTER_REG_17__SCAN_IN) & (P2_INSTADDRPOINTER_REG_18__SCAN_IN | (~new_n1534_ & (new_n1939_ | new_n1940_) & (~new_n1939_ | ~new_n1940_)));
  assign new_n1939_ = (~new_n1330_ | ~P2_EBX_REG_17__SCAN_IN) & new_n1926_ & (~new_n1330_ | ~P2_EBX_REG_15__SCAN_IN) & new_n1924_ & new_n1925_ & (~new_n1330_ | ~P2_EBX_REG_13__SCAN_IN);
  assign new_n1940_ = ~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_18__SCAN_IN);
  assign new_n1941_ = (new_n1942_ | (~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_19__SCAN_IN))) & ~new_n1534_ & (~new_n1942_ | (new_n1330_ & P2_EBX_REG_19__SCAN_IN));
  assign new_n1942_ = new_n1940_ & (~new_n1330_ | ~P2_EBX_REG_17__SCAN_IN) & new_n1926_ & (~new_n1330_ | ~P2_EBX_REG_15__SCAN_IN) & new_n1924_ & new_n1925_ & (~new_n1330_ | ~P2_EBX_REG_13__SCAN_IN);
  assign new_n1943_ = new_n1944_ ^ (new_n1942_ & (~new_n1330_ | ~P2_EBX_REG_19__SCAN_IN));
  assign new_n1944_ = ~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_20__SCAN_IN);
  assign new_n1945_ = ~P2_INSTADDRPOINTER_REG_24__SCAN_IN & (~new_n1946_ | new_n1534_);
  assign new_n1946_ = new_n1949_ ^ (new_n1947_ & (~new_n1330_ | ~P2_EBX_REG_23__SCAN_IN));
  assign new_n1947_ = new_n1948_ & (~new_n1330_ | ~P2_EBX_REG_21__SCAN_IN) & new_n1944_ & new_n1942_ & (~new_n1330_ | ~P2_EBX_REG_19__SCAN_IN);
  assign new_n1948_ = ~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_22__SCAN_IN);
  assign new_n1949_ = ~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_24__SCAN_IN);
  assign new_n1950_ = (~P2_INSTADDRPOINTER_REG_24__SCAN_IN | ~new_n1946_ | new_n1534_) & ((~P2_INSTADDRPOINTER_REG_24__SCAN_IN & (~new_n1946_ | new_n1534_)) | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN | (~new_n1947_ & (new_n1907_ | (new_n1330_ & P2_EBX_REG_23__SCAN_IN))) | new_n1534_ | (new_n1947_ & (~new_n1330_ | ~P2_EBX_REG_23__SCAN_IN)));
  assign new_n1951_ = ((~new_n1941_ & ~P2_INSTADDRPOINTER_REG_19__SCAN_IN) | (~P2_INSTADDRPOINTER_REG_20__SCAN_IN & (~new_n1943_ | new_n1534_)) | ((~new_n1941_ | ~P2_INSTADDRPOINTER_REG_19__SCAN_IN) & (~P2_INSTADDRPOINTER_REG_18__SCAN_IN | new_n1534_ | (new_n1939_ & new_n1940_) | (~new_n1939_ & ~new_n1940_)))) & (~P2_INSTADDRPOINTER_REG_20__SCAN_IN | ~new_n1943_ | new_n1534_);
  assign new_n1952_ = (new_n1954_ | P2_INSTADDRPOINTER_REG_21__SCAN_IN) & (new_n1953_ | P2_INSTADDRPOINTER_REG_22__SCAN_IN);
  assign new_n1953_ = ~new_n1534_ & (~new_n1948_ | (new_n1330_ & P2_EBX_REG_21__SCAN_IN) | ~new_n1944_ | ~new_n1942_ | (new_n1330_ & P2_EBX_REG_19__SCAN_IN)) & (new_n1948_ | ((~new_n1330_ | ~P2_EBX_REG_21__SCAN_IN) & new_n1944_ & new_n1942_ & (~new_n1330_ | ~P2_EBX_REG_19__SCAN_IN)));
  assign new_n1954_ = ~new_n1534_ & (~new_n1330_ | ~P2_EBX_REG_21__SCAN_IN | (~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_20__SCAN_IN) & new_n1942_ & (~new_n1330_ | ~P2_EBX_REG_19__SCAN_IN))) & ~new_n1907_ & ((new_n1330_ & P2_EBX_REG_21__SCAN_IN) | new_n1907_ | (new_n1330_ & P2_EBX_REG_20__SCAN_IN) | ~new_n1942_ | (new_n1330_ & P2_EBX_REG_19__SCAN_IN));
  assign new_n1955_ = (~new_n1953_ | ~P2_INSTADDRPOINTER_REG_22__SCAN_IN) & ((~new_n1953_ & ~P2_INSTADDRPOINTER_REG_22__SCAN_IN) | ~new_n1954_ | ~P2_INSTADDRPOINTER_REG_21__SCAN_IN);
  assign new_n1956_ = ~P2_INSTADDRPOINTER_REG_23__SCAN_IN & ((~new_n1947_ & (new_n1907_ | (new_n1330_ & P2_EBX_REG_23__SCAN_IN))) | new_n1534_ | (new_n1947_ & (~new_n1330_ | ~P2_EBX_REG_23__SCAN_IN)));
  assign new_n1957_ = new_n1974_ & ((~P2_INSTADDRPOINTER_REG_29__SCAN_IN & (~new_n2029_ | ~new_n1958_ | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN)) | ~new_n2028_ | (new_n2029_ & P2_INSTADDRPOINTER_REG_29__SCAN_IN & new_n1958_ & P2_INSTADDRPOINTER_REG_23__SCAN_IN & P2_INSTADDRPOINTER_REG_24__SCAN_IN));
  assign new_n1958_ = new_n1970_ & new_n1959_ & new_n1973_;
  assign new_n1959_ = ((new_n1905_ & P2_INSTADDRPOINTER_REG_8__SCAN_IN) | ((new_n1799_ | P2_INSTADDRPOINTER_REG_7__SCAN_IN) & ((new_n1799_ & P2_INSTADDRPOINTER_REG_7__SCAN_IN) | ((new_n1960_ | P2_INSTADDRPOINTER_REG_6__SCAN_IN) & (new_n1961_ | (new_n1960_ & P2_INSTADDRPOINTER_REG_6__SCAN_IN)))))) & new_n1969_ & (new_n1905_ | P2_INSTADDRPOINTER_REG_8__SCAN_IN);
  assign new_n1960_ = new_n1882_ ^ ~new_n1865_;
  assign new_n1961_ = (new_n1962_ | P2_INSTADDRPOINTER_REG_5__SCAN_IN) & ((new_n1962_ & P2_INSTADDRPOINTER_REG_5__SCAN_IN) | (new_n1963_ & P2_INSTADDRPOINTER_REG_4__SCAN_IN) | ((new_n1963_ | P2_INSTADDRPOINTER_REG_4__SCAN_IN) & ((new_n1964_ & P2_INSTADDRPOINTER_REG_3__SCAN_IN) | (new_n1965_ & (new_n1964_ | P2_INSTADDRPOINTER_REG_3__SCAN_IN)))));
  assign new_n1962_ = ~new_n1860_ ^ (~new_n1855_ & new_n1820_ & new_n1849_);
  assign new_n1963_ = ~new_n1855_ ^ (new_n1820_ & new_n1849_);
  assign new_n1964_ = new_n1820_ ^ new_n1849_;
  assign new_n1965_ = ((P2_INSTADDRPOINTER_REG_2__SCAN_IN & (~new_n1966_ | new_n1967_) & (new_n1966_ | ~new_n1967_)) | (new_n1968_ & P2_INSTADDRPOINTER_REG_1__SCAN_IN) | (new_n1966_ & (~new_n1587_ | ~new_n1322_ | ~new_n1580_) & (new_n1968_ | P2_INSTADDRPOINTER_REG_1__SCAN_IN))) & (P2_INSTADDRPOINTER_REG_2__SCAN_IN | (new_n1966_ ^ ~new_n1967_));
  assign new_n1966_ = ~new_n1848_ & (new_n1322_ | (new_n1821_ & new_n1828_));
  assign new_n1967_ = (~new_n1322_ | new_n1596_) & (~new_n1837_ | ~new_n1841_ | ~new_n1842_);
  assign new_n1968_ = P2_INSTADDRPOINTER_REG_0__SCAN_IN & (new_n1322_ ? new_n1580_ : (~new_n1897_ | ~new_n1898_ | ~new_n1895_ | ~new_n1896_));
  assign new_n1969_ = P2_INSTADDRPOINTER_REG_11__SCAN_IN & P2_INSTADDRPOINTER_REG_12__SCAN_IN & P2_INSTADDRPOINTER_REG_9__SCAN_IN & P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign new_n1970_ = new_n1971_ & new_n1972_;
  assign new_n1971_ = P2_INSTADDRPOINTER_REG_15__SCAN_IN & P2_INSTADDRPOINTER_REG_16__SCAN_IN & P2_INSTADDRPOINTER_REG_17__SCAN_IN & P2_INSTADDRPOINTER_REG_18__SCAN_IN & P2_INSTADDRPOINTER_REG_19__SCAN_IN & P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign new_n1972_ = P2_INSTADDRPOINTER_REG_21__SCAN_IN & P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign new_n1973_ = P2_INSTADDRPOINTER_REG_13__SCAN_IN & P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign new_n1974_ = new_n2014_ & ((new_n2027_ & (~new_n1975_ | ~new_n2023_)) | ~new_n2004_ | (~new_n2027_ & new_n1975_ & new_n2023_));
  assign new_n1975_ = ~new_n2003_ & ~new_n2002_ & ~new_n2001_ & new_n1976_ & ~new_n2000_;
  assign new_n1976_ = ~new_n1999_ & ~new_n1998_ & ~new_n1997_ & ~new_n1996_ & ~new_n1995_ & ~new_n1994_ & new_n1977_ & ~new_n1993_;
  assign new_n1977_ = ~new_n1992_ & ~new_n1991_ & new_n1988_ & ~new_n1987_ & ~new_n1986_ & ~new_n1985_ & new_n1978_ & ~new_n1984_;
  assign new_n1978_ = ~new_n1983_ & ~new_n1982_ & ~new_n1981_ & (new_n1979_ | (~new_n1980_ & (new_n1383_ | (~new_n1386_ & ~new_n1387_))));
  assign new_n1979_ = ((new_n1382_ & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN & (~new_n1328_ | ~new_n1365_))) & (~new_n1379_ | (~new_n1373_ & P2_INSTADDRPOINTER_REG_3__SCAN_IN));
  assign new_n1980_ = (~new_n1382_ | ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | (new_n1328_ & new_n1365_)) & new_n1379_ & (new_n1373_ | ~P2_INSTADDRPOINTER_REG_3__SCAN_IN);
  assign new_n1981_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_4__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_4__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_4__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_4__SCAN_IN);
  assign new_n1982_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_5__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_5__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_5__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_5__SCAN_IN);
  assign new_n1983_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_6__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_6__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_6__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_6__SCAN_IN);
  assign new_n1984_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_7__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_7__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_7__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_7__SCAN_IN);
  assign new_n1985_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_8__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_8__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_8__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_8__SCAN_IN);
  assign new_n1986_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_9__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_9__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_9__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_9__SCAN_IN);
  assign new_n1987_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_10__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_10__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_10__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_10__SCAN_IN);
  assign new_n1988_ = ((~new_n1373_ & P2_INSTADDRPOINTER_REG_11__SCAN_IN) | ~new_n1989_ | (new_n1380_ & P2_REIP_REG_11__SCAN_IN)) & ((~new_n1373_ & P2_INSTADDRPOINTER_REG_12__SCAN_IN) | ~new_n1990_ | (new_n1380_ & P2_REIP_REG_12__SCAN_IN));
  assign new_n1989_ = (~new_n1381_ | ~P2_EBX_REG_11__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_11__SCAN_IN);
  assign new_n1990_ = (~new_n1381_ | ~P2_EBX_REG_12__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_12__SCAN_IN);
  assign new_n1991_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_13__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_13__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_13__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_13__SCAN_IN);
  assign new_n1992_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_14__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_14__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_14__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_14__SCAN_IN);
  assign new_n1993_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_15__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_15__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_15__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_15__SCAN_IN);
  assign new_n1994_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_16__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_16__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_16__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_16__SCAN_IN);
  assign new_n1995_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_17__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_17__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_17__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_17__SCAN_IN);
  assign new_n1996_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_18__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_18__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_18__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_18__SCAN_IN);
  assign new_n1997_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_19__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_19__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_19__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_19__SCAN_IN);
  assign new_n1998_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_20__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_20__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_20__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_20__SCAN_IN);
  assign new_n1999_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_21__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_21__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_21__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_21__SCAN_IN);
  assign new_n2000_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_22__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_22__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_22__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_22__SCAN_IN);
  assign new_n2001_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_23__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_23__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_23__SCAN_IN);
  assign new_n2002_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_24__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_24__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_24__SCAN_IN);
  assign new_n2003_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_25__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_25__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_25__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_25__SCAN_IN);
  assign new_n2004_ = ~new_n2005_ & P2_STATE2_REG_1__SCAN_IN & P2_STATEBS16_REG_SCAN_IN;
  assign new_n2005_ = ~new_n2006_ & ((P2_STATE2_REG_2__SCAN_IN & P2_STATE2_REG_1__SCAN_IN) | P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_0__SCAN_IN);
  assign new_n2006_ = new_n2010_ & (new_n1322_ ? (new_n2009_ & (~new_n1875_ | ~new_n1782_ | ~new_n2007_ | new_n2008_)) : new_n2011_);
  assign new_n2007_ = new_n1764_ ? ~new_n1607_ : new_n1779_;
  assign new_n2008_ = ((new_n1587_ & new_n1764_) | (~new_n1764_ & ~new_n1772_) | (~new_n1764_ & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (new_n1764_ ? new_n1580_ : (~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))) & (new_n1764_ ? new_n1596_ : new_n1774_);
  assign new_n2009_ = (~new_n1551_ | ~new_n1764_) ^ ((~new_n1560_ | ~new_n1764_) & ((~new_n1764_ & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) | (((~new_n1764_ & new_n1765_) | (~new_n1764_ & new_n1766_)) & (new_n1764_ ? ~new_n1569_ : (P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)))));
  assign new_n2010_ = new_n1791_ & ~new_n1370_ & new_n1356_ & new_n1367_ & ~new_n1317_ & ~new_n1330_ & new_n1350_;
  assign new_n2011_ = ((~new_n2012_ & P2_STATE2_REG_1__SCAN_IN) | ((~new_n2013_ | ~new_n1779_ | (new_n1767_ ^ (~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ^ ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN))) & ~P2_STATE2_REG_1__SCAN_IN & ((~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) | (~new_n1767_ & (~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN))))) & (P2_FLUSH_REG_SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  assign new_n2012_ = (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & ~P2_FLUSH_REG_SCAN_IN & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign new_n2013_ = ((P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) ^ ((~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | ((~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)))) & ((~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) ? (~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) : (P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN));
  assign new_n2014_ = ((~new_n2015_ & ~P2_PHYADDRPOINTER_REG_29__SCAN_IN) | new_n2005_ | new_n2021_ | (new_n2015_ & P2_PHYADDRPOINTER_REG_29__SCAN_IN)) & (~new_n2005_ | ~P2_PHYADDRPOINTER_REG_29__SCAN_IN) & (~P2_REIP_REG_29__SCAN_IN | new_n2005_ | ~new_n2022_);
  assign new_n2015_ = P2_PHYADDRPOINTER_REG_28__SCAN_IN & P2_PHYADDRPOINTER_REG_26__SCAN_IN & P2_PHYADDRPOINTER_REG_27__SCAN_IN & new_n2016_ & P2_PHYADDRPOINTER_REG_25__SCAN_IN;
  assign new_n2016_ = new_n2017_ & P2_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign new_n2017_ = P2_PHYADDRPOINTER_REG_23__SCAN_IN & P2_PHYADDRPOINTER_REG_22__SCAN_IN & P2_PHYADDRPOINTER_REG_21__SCAN_IN & P2_PHYADDRPOINTER_REG_20__SCAN_IN & P2_PHYADDRPOINTER_REG_19__SCAN_IN & P2_PHYADDRPOINTER_REG_18__SCAN_IN & new_n2018_ & P2_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign new_n2018_ = P2_PHYADDRPOINTER_REG_16__SCAN_IN & P2_PHYADDRPOINTER_REG_15__SCAN_IN & P2_PHYADDRPOINTER_REG_14__SCAN_IN & P2_PHYADDRPOINTER_REG_13__SCAN_IN & new_n2020_ & P2_PHYADDRPOINTER_REG_10__SCAN_IN & new_n2019_ & P2_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign new_n2019_ = P2_PHYADDRPOINTER_REG_8__SCAN_IN & P2_PHYADDRPOINTER_REG_7__SCAN_IN & P2_PHYADDRPOINTER_REG_6__SCAN_IN & P2_PHYADDRPOINTER_REG_5__SCAN_IN & P2_PHYADDRPOINTER_REG_4__SCAN_IN & P2_PHYADDRPOINTER_REG_3__SCAN_IN & P2_PHYADDRPOINTER_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign new_n2020_ = P2_PHYADDRPOINTER_REG_11__SCAN_IN & P2_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign new_n2021_ = ~new_n1407_ & (~P2_STATE2_REG_1__SCAN_IN | P2_STATEBS16_REG_SCAN_IN);
  assign new_n2022_ = ~P2_STATE2_REG_2__SCAN_IN & ~P2_STATE2_REG_1__SCAN_IN;
  assign new_n2023_ = (~new_n2024_ | (~new_n1373_ & P2_INSTADDRPOINTER_REG_28__SCAN_IN)) & (~new_n2026_ | (~new_n1373_ & P2_INSTADDRPOINTER_REG_27__SCAN_IN)) & (~new_n2025_ | (~new_n1373_ & P2_INSTADDRPOINTER_REG_26__SCAN_IN));
  assign new_n2024_ = (~new_n1381_ | ~P2_EBX_REG_28__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_28__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_28__SCAN_IN);
  assign new_n2025_ = (~new_n1380_ | ~P2_REIP_REG_26__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_26__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_26__SCAN_IN);
  assign new_n2026_ = (~new_n1380_ | ~P2_REIP_REG_27__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_27__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_27__SCAN_IN);
  assign new_n2027_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_29__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_29__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_29__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_29__SCAN_IN);
  assign new_n2028_ = ~new_n2005_ & new_n1322_ & P2_STATE2_REG_0__SCAN_IN;
  assign new_n2029_ = P2_INSTADDRPOINTER_REG_27__SCAN_IN & P2_INSTADDRPOINTER_REG_28__SCAN_IN & P2_INSTADDRPOINTER_REG_25__SCAN_IN & P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign new_n2030_ = new_n2031_ ^ P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign new_n2031_ = (new_n2032_ | (~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_29__SCAN_IN))) & ~new_n1534_ & (~new_n2032_ | (new_n1330_ & P2_EBX_REG_29__SCAN_IN));
  assign new_n2032_ = ~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_28__SCAN_IN) & (~new_n1330_ | ~P2_EBX_REG_27__SCAN_IN) & new_n2033_ & (~new_n1330_ | ~P2_EBX_REG_25__SCAN_IN) & (~new_n1330_ | ~P2_EBX_REG_26__SCAN_IN);
  assign new_n2033_ = new_n1949_ & (~new_n1330_ | ~P2_EBX_REG_23__SCAN_IN) & new_n1948_ & (~new_n1330_ | ~P2_EBX_REG_21__SCAN_IN) & new_n1944_ & new_n1942_ & (~new_n1330_ | ~P2_EBX_REG_19__SCAN_IN);
  assign new_n2034_ = (new_n2035_ | P2_INSTADDRPOINTER_REG_28__SCAN_IN) & (new_n2037_ | P2_INSTADDRPOINTER_REG_26__SCAN_IN) & (new_n2036_ | P2_INSTADDRPOINTER_REG_27__SCAN_IN);
  assign new_n2035_ = (((~new_n1330_ | ~P2_EBX_REG_27__SCAN_IN) & ~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_26__SCAN_IN) & new_n2033_ & (~new_n1330_ | ~P2_EBX_REG_25__SCAN_IN)) | (~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_28__SCAN_IN))) & ~new_n1534_ & ((new_n1330_ & P2_EBX_REG_27__SCAN_IN) | new_n1907_ | (new_n1330_ & P2_EBX_REG_26__SCAN_IN) | ~new_n2033_ | (new_n1330_ & P2_EBX_REG_25__SCAN_IN) | (new_n1330_ & P2_EBX_REG_28__SCAN_IN));
  assign new_n2036_ = ((~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_26__SCAN_IN) & new_n2033_ & (~new_n1330_ | ~P2_EBX_REG_25__SCAN_IN)) | (~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_27__SCAN_IN))) & ~new_n1534_ & ((new_n1330_ & P2_EBX_REG_27__SCAN_IN) | new_n1907_ | (new_n1330_ & P2_EBX_REG_26__SCAN_IN) | ~new_n2033_ | (new_n1330_ & P2_EBX_REG_25__SCAN_IN));
  assign new_n2037_ = ((~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_26__SCAN_IN)) | (new_n2033_ & (~new_n1330_ | ~P2_EBX_REG_25__SCAN_IN))) & ~new_n1534_ & (new_n1907_ | (new_n1330_ & P2_EBX_REG_26__SCAN_IN) | ~new_n2033_ | (new_n1330_ & P2_EBX_REG_25__SCAN_IN));
  assign new_n2038_ = (~new_n2035_ | ~P2_INSTADDRPOINTER_REG_28__SCAN_IN) & ((~new_n2035_ & ~P2_INSTADDRPOINTER_REG_28__SCAN_IN) | ((~new_n2036_ | ~P2_INSTADDRPOINTER_REG_27__SCAN_IN) & (~new_n2037_ | ~P2_INSTADDRPOINTER_REG_26__SCAN_IN | (~new_n2036_ & ~P2_INSTADDRPOINTER_REG_27__SCAN_IN))));
  assign new_n2039_ = ~new_n1534_ & (new_n2033_ | ~new_n1330_ | ~P2_EBX_REG_25__SCAN_IN) & ~new_n1907_ & (~new_n2033_ | (new_n1330_ & P2_EBX_REG_25__SCAN_IN));
  assign new_n2040_ = ~new_n2005_ & ~new_n1322_ & P2_STATE2_REG_0__SCAN_IN;
  assign new_n2041_ = (new_n2042_ | ~new_n2476_ | new_n2053_) & (new_n2476_ | ~P1_EBX_REG_29__SCAN_IN) & ((~new_n2498_ & (~new_n2450_ | ~new_n2496_)) | ~new_n2476_ | ~new_n2053_ | (new_n2498_ & new_n2450_ & new_n2496_));
  assign new_n2042_ = ~new_n2439_ ^ (~new_n2043_ & ~new_n2449_);
  assign new_n2043_ = (((~new_n2324_ | ~new_n2425_) & ((~new_n2324_ & ~new_n2425_) | ((~new_n2324_ | ~new_n2432_) & ((~new_n2044_ & new_n2422_) | (~new_n2324_ & ~new_n2432_))))) | ~new_n2423_ | (~new_n2324_ & ~new_n2424_)) & (new_n2367_ | (~new_n2324_ & ~new_n2424_));
  assign new_n2044_ = ((new_n2324_ & new_n2346_) | ((new_n2324_ | new_n2346_) & ((new_n2324_ & ~new_n2339_) | ((new_n2324_ | ~new_n2339_) & (new_n2327_ | (~new_n2045_ & ~new_n2338_)))))) & (new_n2324_ | new_n2360_) & (new_n2324_ | ~new_n2353_);
  assign new_n2045_ = new_n2323_ & (~new_n2308_ | (~new_n2046_ & (new_n2242_ | (~new_n2243_ & (new_n2248_ | (~new_n2249_ & new_n2304_))))));
  assign new_n2046_ = ~new_n2239_ & new_n2237_ & ((new_n2227_ ^ ~new_n2163_) | ~new_n2047_ | (~new_n2232_ ^ new_n2163_)) & ((new_n2227_ & ~new_n2163_) | (~new_n2227_ & new_n2163_) | (new_n2047_ & (new_n2232_ ^ new_n2163_)));
  assign new_n2047_ = ~new_n2202_ & ~new_n2209_ & ~new_n2215_ & ~new_n2048_ & ~new_n2221_;
  assign new_n2048_ = new_n2191_ & (~new_n2177_ | new_n2201_ | (~new_n2049_ & (new_n2147_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_))))));
  assign new_n2049_ = ~new_n2135_ & (new_n2145_ | (~P1_STATE2_REG_0__SCAN_IN & (new_n2133_ | new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_)))) & (~new_n2133_ | (~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))))));
  assign new_n2050_ = new_n2117_ & (~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (new_n2051_ & new_n2105_ & new_n2110_));
  assign new_n2051_ = (~P1_STATE2_REG_0__SCAN_IN | (~new_n2052_ & (new_n2097_ | (~new_n2090_ & new_n2073_)))) & (~new_n2096_ | ~P1_STATE2_REG_0__SCAN_IN) & (new_n2104_ | ~new_n2090_ | new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN);
  assign new_n2052_ = new_n2067_ & ~new_n2073_ & (new_n2053_ | (new_n2065_ & ~new_n2085_) | ~new_n2079_ | (~new_n2060_ & new_n2085_));
  assign new_n2053_ = new_n2054_ & new_n2058_ & new_n2059_ & new_n2055_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_15__7__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_11__7__SCAN_IN);
  assign new_n2054_ = (~P1_INSTQUEUE_REG_6__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P1_INSTQUEUE_REG_7__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2055_ = (~P1_INSTQUEUE_REG_9__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_4__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_2__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2056_ = P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign new_n2057_ = P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign new_n2058_ = (~P1_INSTQUEUE_REG_1__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_8__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_5__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2059_ = (~P1_INSTQUEUE_REG_14__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_0__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2060_ = new_n2061_ & new_n2062_ & new_n2063_ & new_n2064_;
  assign new_n2061_ = (~P1_INSTQUEUE_REG_15__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_6__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P1_INSTQUEUE_REG_11__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2062_ = (~P1_INSTQUEUE_REG_8__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_4__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_5__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2063_ = (~P1_INSTQUEUE_REG_1__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_2__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2064_ = (~P1_INSTQUEUE_REG_3__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_9__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_10__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2065_ = (~new_n2066_ | ~P1_INSTQUEUE_REG_0__5__SCAN_IN) & new_n2061_ & new_n2062_ & new_n2063_ & new_n2064_;
  assign new_n2066_ = ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign new_n2067_ = new_n2068_ & new_n2071_ & new_n2072_ & new_n2069_ & new_n2070_;
  assign new_n2068_ = (~P1_INSTQUEUE_REG_15__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2069_ = (~P1_INSTQUEUE_REG_10__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_5__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_1__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_14__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2070_ = (~P1_INSTQUEUE_REG_3__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_6__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2071_ = (~P1_INSTQUEUE_REG_9__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_4__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_2__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2072_ = (~P1_INSTQUEUE_REG_8__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_12__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_0__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2073_ = new_n2074_ & new_n2077_ & new_n2078_ & new_n2075_ & new_n2076_;
  assign new_n2074_ = (~P1_INSTQUEUE_REG_6__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P1_INSTQUEUE_REG_7__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2075_ = (~P1_INSTQUEUE_REG_2__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_9__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_12__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_4__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2076_ = (~P1_INSTQUEUE_REG_15__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2077_ = (~P1_INSTQUEUE_REG_5__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_8__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_10__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2078_ = (~P1_INSTQUEUE_REG_14__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_1__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_0__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2079_ = new_n2081_ & new_n2083_ & new_n2084_ & new_n2082_ & (~new_n2080_ | ~P1_INSTQUEUE_REG_7__4__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_11__4__SCAN_IN);
  assign new_n2080_ = ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign new_n2081_ = (~P1_INSTQUEUE_REG_6__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P1_INSTQUEUE_REG_3__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_15__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2082_ = (P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ((~P1_INSTQUEUE_REG_0__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_8__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN))) & (~P1_INSTQUEUE_REG_4__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2083_ = (~P1_INSTQUEUE_REG_2__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2084_ = (~P1_INSTQUEUE_REG_9__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_1__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_5__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2085_ = new_n2086_ & ~new_n2088_ & new_n2089_ & new_n2087_ & (~new_n2080_ | ~P1_INSTQUEUE_REG_7__6__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_11__6__SCAN_IN);
  assign new_n2086_ = (~P1_INSTQUEUE_REG_3__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_6__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P1_INSTQUEUE_REG_15__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2087_ = (~P1_INSTQUEUE_REG_14__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_1__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_9__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2088_ = ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ((P1_INSTQUEUE_REG_0__6__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (P1_INSTQUEUE_REG_8__6__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | (P1_INSTQUEUE_REG_12__6__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n2089_ = (~P1_INSTQUEUE_REG_5__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_10__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_4__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_2__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2090_ = ~new_n2067_ & ~new_n2091_;
  assign new_n2091_ = new_n2092_ & new_n2094_ & new_n2095_ & new_n2093_ & (~new_n2057_ | ~P1_INSTQUEUE_REG_11__3__SCAN_IN) & (~new_n2056_ | ~P1_INSTQUEUE_REG_15__3__SCAN_IN);
  assign new_n2092_ = (~P1_INSTQUEUE_REG_6__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P1_INSTQUEUE_REG_7__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2093_ = (~P1_INSTQUEUE_REG_9__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_4__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_2__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2094_ = (~P1_INSTQUEUE_REG_1__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_8__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_5__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2095_ = (~P1_INSTQUEUE_REG_14__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_0__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2096_ = ~new_n2053_ & ~new_n2085_ & new_n2097_ & new_n2091_ & new_n2065_ & new_n2067_ & new_n2073_;
  assign new_n2097_ = new_n2100_ & new_n2102_ & new_n2103_ & new_n2101_ & (~new_n2098_ | ~P1_INSTQUEUE_REG_6__2__SCAN_IN) & (~new_n2099_ | ~P1_INSTQUEUE_REG_3__2__SCAN_IN);
  assign new_n2098_ = ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign new_n2099_ = ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign new_n2100_ = (~P1_INSTQUEUE_REG_15__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2101_ = (~P1_INSTQUEUE_REG_2__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_1__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_5__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2102_ = (~P1_INSTQUEUE_REG_13__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_4__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_9__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2103_ = (~P1_INSTQUEUE_REG_8__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_0__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2104_ = (new_n2079_ | (~new_n2065_ & new_n2085_)) & ~new_n2053_ & (~new_n2065_ | new_n2085_) & (~new_n2085_ | new_n2065_ | ~new_n2079_);
  assign new_n2105_ = (~new_n2107_ | ~P1_STATE2_REG_0__SCAN_IN) & (~new_n2106_ | ~new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN) & new_n2109_ & (~new_n2108_ | ~P1_STATE2_REG_0__SCAN_IN);
  assign new_n2106_ = new_n2097_ & new_n2091_ & ~new_n2085_ & new_n2065_ & new_n2053_ & new_n2079_;
  assign new_n2107_ = ~new_n2067_ & ~new_n2091_ & ~new_n2053_ & ~new_n2085_ & ~new_n2065_ & new_n2079_;
  assign new_n2108_ = ~new_n2097_ & new_n2085_ & new_n2065_ & new_n2053_ & new_n2079_;
  assign new_n2109_ = (~P1_STATE2_REG_0__SCAN_IN | new_n2067_ | ~new_n2073_) & (~new_n2091_ | new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN);
  assign new_n2110_ = (~new_n2111_ | ((new_n2097_ | ((~new_n2065_ | new_n2085_) & new_n2079_ & (new_n2053_ | ~new_n2085_))) & (new_n2097_ | ~new_n2091_ | new_n2065_ | ~new_n2079_ | new_n2053_ | new_n2085_) & (~new_n2097_ | ~new_n2091_ | new_n2053_ | new_n2079_ | ~new_n2085_))) & ~new_n2113_ & (~new_n2111_ | ((new_n2091_ | (~new_n2065_ & ~new_n2053_ & ~new_n2079_ & new_n2085_)) & (~new_n2053_ | (new_n2065_ & new_n2079_)) & ((new_n2065_ & ~new_n2085_) | ~new_n2097_ | (~new_n2079_ & new_n2085_))));
  assign new_n2111_ = new_n2073_ & new_n2112_;
  assign new_n2112_ = P1_STATE2_REG_0__SCAN_IN & new_n2068_ & new_n2071_ & new_n2072_ & new_n2069_ & new_n2070_;
  assign new_n2113_ = new_n2114_ & ~new_n2115_ & new_n2065_ & new_n2079_ & ~new_n2053_ & new_n2085_ & new_n2097_ & ~new_n2091_;
  assign new_n2114_ = P1_STATE2_REG_0__SCAN_IN & (~new_n2074_ | ~new_n2077_ | ~new_n2078_ | ~new_n2075_ | ~new_n2076_);
  assign new_n2115_ = new_n2116_ & new_n2068_ & new_n2071_ & new_n2072_ & new_n2069_ & new_n2070_;
  assign new_n2116_ = P1_STATE_REG_2__SCAN_IN ^ ~P1_STATE_REG_1__SCAN_IN;
  assign new_n2117_ = (new_n2118_ | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~new_n2119_ | ~new_n2120_);
  assign new_n2118_ = P1_STATE2_REG_2__SCAN_IN & ~P1_STATE2_REG_1__SCAN_IN;
  assign new_n2119_ = ~P1_STATE2_REG_0__SCAN_IN & ~P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_1__SCAN_IN;
  assign new_n2120_ = P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ^ P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n2121_ = ~new_n2122_ & (new_n2130_ | (P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & (new_n2127_ | ~new_n2051_ | ~new_n2128_)));
  assign new_n2122_ = ~new_n2123_ & ~new_n2124_ & ~new_n2125_ & ~new_n2107_ & new_n2126_ & (~new_n2108_ | ~new_n2091_);
  assign new_n2123_ = (~new_n2067_ | (~new_n2091_ & (new_n2065_ | new_n2053_ | new_n2079_ | ~new_n2085_)) | (new_n2053_ & (~new_n2065_ | ~new_n2079_)) | ((~new_n2065_ | new_n2085_) & new_n2097_ & (new_n2079_ | ~new_n2085_)) | (~new_n2097_ & ((new_n2065_ & ~new_n2085_) | ~new_n2079_ | (~new_n2053_ & new_n2085_)))) & new_n2073_ & (~new_n2079_ | new_n2065_ | new_n2067_);
  assign new_n2124_ = (~new_n2067_ | (~new_n2073_ & (~new_n2079_ | new_n2091_ | (new_n2065_ & ~new_n2085_) | ((new_n2053_ | ~new_n2065_) & (new_n2053_ | new_n2085_))))) & ((~new_n2079_ & (new_n2065_ | ~new_n2085_)) | new_n2053_ | (new_n2065_ & ~new_n2085_) | (new_n2085_ & ~new_n2065_ & new_n2079_) | new_n2067_ | new_n2073_ | (new_n2097_ & new_n2091_));
  assign new_n2125_ = new_n2073_ & new_n2097_ & new_n2091_ & ((~new_n2053_ & ~new_n2079_ & new_n2085_) | (~new_n2085_ & new_n2065_ & new_n2053_ & new_n2079_));
  assign new_n2126_ = (new_n2073_ | new_n2097_) & P1_STATE2_REG_0__SCAN_IN & ~P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_1__SCAN_IN;
  assign new_n2127_ = new_n2111_ & ((new_n2097_ & new_n2091_ & ~new_n2053_ & ~new_n2079_ & new_n2085_) | (~new_n2091_ & (new_n2065_ | new_n2053_ | new_n2079_ | ~new_n2085_)) | (new_n2053_ & (~new_n2065_ | ~new_n2079_)) | ((~new_n2065_ | new_n2085_) & new_n2097_ & (new_n2079_ | ~new_n2085_)) | (~new_n2097_ & ((new_n2065_ & ~new_n2085_) | ~new_n2079_ | (~new_n2053_ & new_n2085_))));
  assign new_n2128_ = ~new_n2113_ & ~new_n2129_ & (~new_n2107_ | ~P1_STATE2_REG_0__SCAN_IN) & new_n2109_ & (~new_n2108_ | ~P1_STATE2_REG_0__SCAN_IN) & (~new_n2106_ | ~new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN);
  assign new_n2129_ = new_n2073_ & new_n2112_ & ~new_n2097_ & new_n2091_ & ~new_n2053_ & ~new_n2085_ & ~new_n2065_ & new_n2079_;
  assign new_n2130_ = P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ? ~new_n2118_ : new_n2119_;
  assign new_n2131_ = new_n2132_ & (~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | (~new_n2127_ & new_n2051_ & new_n2128_));
  assign new_n2132_ = (new_n2118_ | ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (~new_n2119_ | (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)));
  assign new_n2133_ = new_n2134_ & (~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | (~new_n2127_ & new_n2051_ & new_n2128_));
  assign new_n2134_ = (new_n2118_ | ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) & (~new_n2119_ | (P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ^ (~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)));
  assign new_n2135_ = (~new_n2137_ | new_n2138_) & (~new_n2136_ | ~P1_INSTQUEUE_REG_0__3__SCAN_IN);
  assign new_n2136_ = new_n2114_ & ~new_n2079_;
  assign new_n2137_ = new_n2073_ & P1_STATE2_REG_0__SCAN_IN;
  assign new_n2138_ = new_n2139_ & new_n2140_ & new_n2142_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_0__3__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_7__3__SCAN_IN);
  assign new_n2139_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_4__3__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_12__3__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_8__3__SCAN_IN);
  assign new_n2140_ = new_n2141_ & (~P1_INSTQUEUE_REG_9__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_3__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2141_ = (~P1_INSTQUEUE_REG_5__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_15__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_1__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2142_ = (~P1_INSTQUEUE_REG_6__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_2__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2143_ = ~new_n2113_ & ~new_n2129_ & (~new_n2144_ | ~new_n2073_ | ~new_n2097_ | ~new_n2091_);
  assign new_n2144_ = new_n2065_ & P1_STATE2_REG_0__SCAN_IN & new_n2067_ & ~new_n2053_ & ~new_n2085_;
  assign new_n2145_ = new_n2146_ & ~new_n2138_;
  assign new_n2146_ = new_n2079_ & P1_STATE2_REG_0__SCAN_IN;
  assign new_n2147_ = new_n2135_ & ~new_n2145_ & (P1_STATE2_REG_0__SCAN_IN | (~new_n2133_ & ~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))) | (new_n2133_ & (new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_))))));
  assign new_n2148_ = (P1_STATE2_REG_0__SCAN_IN | (~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))) | (new_n2131_ & (new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_)))) & (new_n2149_ | ~new_n2079_ | ~P1_STATE2_REG_0__SCAN_IN);
  assign new_n2149_ = new_n2150_ & new_n2151_ & new_n2153_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_0__2__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_7__2__SCAN_IN);
  assign new_n2150_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_4__2__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_12__2__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_8__2__SCAN_IN);
  assign new_n2151_ = new_n2152_ & (~P1_INSTQUEUE_REG_9__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_3__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2152_ = (~P1_INSTQUEUE_REG_5__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_15__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_1__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2153_ = (~P1_INSTQUEUE_REG_6__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_2__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2154_ = (new_n2175_ | (~new_n2169_ & (P1_STATE2_REG_0__SCAN_IN | (new_n2121_ ^ ~new_n2155_)))) & ((~new_n2163_ & (new_n2156_ | new_n2176_)) | (new_n2175_ & ~new_n2169_ & (P1_STATE2_REG_0__SCAN_IN | (new_n2121_ ^ ~new_n2155_))));
  assign new_n2155_ = ~new_n2143_ ^ (~new_n2117_ | (P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & (~new_n2051_ | ~new_n2105_ | ~new_n2110_)));
  assign new_n2156_ = ~new_n2157_ & (P1_STATE2_REG_0__SCAN_IN | (~new_n2122_ & (new_n2130_ | (P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & (new_n2127_ | ~new_n2051_ | ~new_n2128_)))) | (new_n2122_ & ~new_n2130_ & (~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~new_n2127_ & new_n2051_ & new_n2128_))));
  assign new_n2157_ = new_n2146_ & ~new_n2158_;
  assign new_n2158_ = new_n2159_ & new_n2160_ & new_n2162_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_0__0__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_7__0__SCAN_IN);
  assign new_n2159_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_4__0__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_8__0__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_12__0__SCAN_IN);
  assign new_n2160_ = new_n2161_ & (~P1_INSTQUEUE_REG_9__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_3__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2161_ = (~P1_INSTQUEUE_REG_5__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_15__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_1__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2162_ = (~P1_INSTQUEUE_REG_6__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_2__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2163_ = new_n2146_ & ~new_n2164_;
  assign new_n2164_ = new_n2165_ & new_n2166_ & new_n2168_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_0__7__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_7__7__SCAN_IN);
  assign new_n2165_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_4__7__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_12__7__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_8__7__SCAN_IN);
  assign new_n2166_ = new_n2167_ & (~P1_INSTQUEUE_REG_9__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_3__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2167_ = (~P1_INSTQUEUE_REG_5__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_15__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_1__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2168_ = (~P1_INSTQUEUE_REG_6__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_2__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2169_ = new_n2146_ & ~new_n2170_;
  assign new_n2170_ = new_n2171_ & new_n2172_ & new_n2174_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_0__1__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_7__1__SCAN_IN);
  assign new_n2171_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_4__1__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_12__1__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_8__1__SCAN_IN);
  assign new_n2172_ = new_n2173_ & (~P1_INSTQUEUE_REG_9__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_3__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2173_ = (~P1_INSTQUEUE_REG_5__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_15__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_1__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2174_ = (~P1_INSTQUEUE_REG_6__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_2__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2175_ = (~P1_INSTQUEUE_REG_0__1__SCAN_IN | new_n2079_ | new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN) & (~new_n2164_ | ~new_n2079_ | ~P1_STATE2_REG_0__SCAN_IN) & (new_n2170_ | ~new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN);
  assign new_n2176_ = (~P1_INSTQUEUE_REG_0__0__SCAN_IN | new_n2073_ | new_n2079_) & (new_n2158_ | ~new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN) & P1_STATE2_REG_0__SCAN_IN & (new_n2164_ | ~new_n2079_);
  assign new_n2177_ = ~new_n2185_ & ~new_n2178_ & (new_n2163_ | ~new_n2184_);
  assign new_n2178_ = (~P1_INSTQUEUE_REG_0__6__SCAN_IN | new_n2079_ | new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN) & (new_n2179_ | ~new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN) & (new_n2179_ | ~new_n2079_ | ~P1_STATE2_REG_0__SCAN_IN);
  assign new_n2179_ = new_n2180_ & new_n2181_ & new_n2183_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_0__6__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_7__6__SCAN_IN);
  assign new_n2180_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_4__6__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_12__6__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_8__6__SCAN_IN);
  assign new_n2181_ = new_n2182_ & (~P1_INSTQUEUE_REG_9__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_3__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2182_ = (~P1_INSTQUEUE_REG_5__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_15__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_1__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2183_ = (~P1_INSTQUEUE_REG_6__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_2__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2184_ = (new_n2164_ | ~new_n2137_) & (~new_n2136_ | ~P1_INSTQUEUE_REG_0__7__SCAN_IN);
  assign new_n2185_ = (~P1_INSTQUEUE_REG_0__5__SCAN_IN | new_n2079_ | new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN) & (new_n2186_ | ~new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN) & (new_n2186_ | ~new_n2079_ | ~P1_STATE2_REG_0__SCAN_IN);
  assign new_n2186_ = new_n2187_ & new_n2188_ & new_n2190_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_0__5__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_7__5__SCAN_IN);
  assign new_n2187_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_4__5__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_12__5__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_8__5__SCAN_IN);
  assign new_n2188_ = new_n2189_ & (~P1_INSTQUEUE_REG_9__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_3__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2189_ = (~P1_INSTQUEUE_REG_5__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_15__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_1__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2190_ = (~P1_INSTQUEUE_REG_6__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_2__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2191_ = (~new_n2163_ | new_n2184_) & (new_n2178_ | (~new_n2163_ & new_n2184_) | (~new_n2198_ & ~new_n2199_ & (new_n2185_ | ~new_n2192_)));
  assign new_n2192_ = ((P1_INSTQUEUE_REG_0__4__SCAN_IN & ~new_n2079_ & ~new_n2073_ & P1_STATE2_REG_0__SCAN_IN) | (~new_n2193_ & new_n2073_ & P1_STATE2_REG_0__SCAN_IN)) & ~new_n2193_ & new_n2079_ & P1_STATE2_REG_0__SCAN_IN;
  assign new_n2193_ = new_n2194_ & new_n2195_ & new_n2197_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_0__4__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_7__4__SCAN_IN);
  assign new_n2194_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_4__4__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_12__4__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_8__4__SCAN_IN);
  assign new_n2195_ = new_n2196_ & (~P1_INSTQUEUE_REG_9__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_3__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2196_ = (~P1_INSTQUEUE_REG_5__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_15__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_1__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2197_ = (~P1_INSTQUEUE_REG_6__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_2__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2198_ = ((P1_INSTQUEUE_REG_0__5__SCAN_IN & ~new_n2079_ & ~new_n2073_ & P1_STATE2_REG_0__SCAN_IN) | (~new_n2186_ & new_n2073_ & P1_STATE2_REG_0__SCAN_IN)) & ~new_n2186_ & new_n2079_ & P1_STATE2_REG_0__SCAN_IN;
  assign new_n2199_ = ((P1_INSTQUEUE_REG_0__6__SCAN_IN & ~new_n2079_ & ~new_n2073_ & P1_STATE2_REG_0__SCAN_IN) | (~new_n2179_ & new_n2073_ & P1_STATE2_REG_0__SCAN_IN)) & ~new_n2179_ & new_n2079_ & P1_STATE2_REG_0__SCAN_IN;
  assign new_n2200_ = (~new_n2137_ | new_n2149_) & (~new_n2136_ | ~P1_INSTQUEUE_REG_0__2__SCAN_IN);
  assign new_n2201_ = (~P1_INSTQUEUE_REG_0__4__SCAN_IN | new_n2079_ | new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN) & (new_n2193_ | ~new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN) & (new_n2193_ | ~new_n2079_ | ~P1_STATE2_REG_0__SCAN_IN);
  assign new_n2202_ = new_n2203_ ^ ~new_n2163_;
  assign new_n2203_ = ~new_n2204_ & (~new_n2205_ | ~new_n2206_ | ~new_n2208_ | (new_n2056_ & P1_INSTQUEUE_REG_1__3__SCAN_IN) | (new_n2080_ & P1_INSTQUEUE_REG_9__3__SCAN_IN));
  assign new_n2204_ = ~new_n2136_ & ~new_n2137_;
  assign new_n2205_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_5__3__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_13__3__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_8__3__SCAN_IN);
  assign new_n2206_ = new_n2207_ & (~P1_INSTQUEUE_REG_15__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_6__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2207_ = (~P1_INSTQUEUE_REG_4__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_0__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2208_ = (~P1_INSTQUEUE_REG_2__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_14__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2209_ = new_n2210_ ^ ~new_n2163_;
  assign new_n2210_ = ~new_n2204_ & (~new_n2211_ | ~new_n2212_ | ~new_n2214_ | (new_n2056_ & P1_INSTQUEUE_REG_1__2__SCAN_IN) | (new_n2080_ & P1_INSTQUEUE_REG_9__2__SCAN_IN));
  assign new_n2211_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_5__2__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_13__2__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_8__2__SCAN_IN);
  assign new_n2212_ = new_n2213_ & (~P1_INSTQUEUE_REG_15__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_6__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2213_ = (~P1_INSTQUEUE_REG_4__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_0__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2214_ = (~P1_INSTQUEUE_REG_2__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_14__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2215_ = new_n2216_ ^ ~new_n2163_;
  assign new_n2216_ = ~new_n2204_ & (~new_n2217_ | ~new_n2218_ | ~new_n2220_ | (new_n2056_ & P1_INSTQUEUE_REG_1__1__SCAN_IN) | (new_n2080_ & P1_INSTQUEUE_REG_9__1__SCAN_IN));
  assign new_n2217_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_5__1__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_13__1__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_8__1__SCAN_IN);
  assign new_n2218_ = new_n2219_ & (~P1_INSTQUEUE_REG_15__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_6__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2219_ = (~P1_INSTQUEUE_REG_4__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_0__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2220_ = (~P1_INSTQUEUE_REG_2__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_14__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2221_ = new_n2222_ ^ ~new_n2163_;
  assign new_n2222_ = ~new_n2204_ & (~new_n2223_ | ~new_n2224_ | ~new_n2226_ | (new_n2056_ & P1_INSTQUEUE_REG_1__0__SCAN_IN) | (new_n2080_ & P1_INSTQUEUE_REG_9__0__SCAN_IN));
  assign new_n2223_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_5__0__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_13__0__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_8__0__SCAN_IN);
  assign new_n2224_ = new_n2225_ & (~P1_INSTQUEUE_REG_15__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_6__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2225_ = (~P1_INSTQUEUE_REG_4__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_11__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_0__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2226_ = (~P1_INSTQUEUE_REG_2__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_14__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2227_ = ~new_n2204_ & (~new_n2228_ | ~new_n2229_ | ~new_n2231_ | (new_n2056_ & P1_INSTQUEUE_REG_1__5__SCAN_IN) | (new_n2080_ & P1_INSTQUEUE_REG_9__5__SCAN_IN));
  assign new_n2228_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_5__5__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_13__5__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_8__5__SCAN_IN);
  assign new_n2229_ = new_n2230_ & (~P1_INSTQUEUE_REG_15__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_6__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2230_ = (~P1_INSTQUEUE_REG_4__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_0__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2231_ = (~P1_INSTQUEUE_REG_2__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_14__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2232_ = ~new_n2204_ & (~new_n2233_ | ~new_n2234_ | ~new_n2236_ | (new_n2056_ & P1_INSTQUEUE_REG_1__4__SCAN_IN) | (new_n2080_ & P1_INSTQUEUE_REG_9__4__SCAN_IN));
  assign new_n2233_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_5__4__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_13__4__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_8__4__SCAN_IN);
  assign new_n2234_ = new_n2235_ & (~P1_INSTQUEUE_REG_15__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_6__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2235_ = (~P1_INSTQUEUE_REG_4__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_0__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2236_ = (~P1_INSTQUEUE_REG_2__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_14__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2237_ = ~new_n2238_ & P1_STATE2_REG_2__SCAN_IN;
  assign new_n2238_ = new_n2067_ & ~new_n2085_;
  assign new_n2239_ = (~P1_EAX_REG_13__SCAN_IN | ~new_n2053_ | ~P1_STATE2_REG_2__SCAN_IN) & ((P1_PHYADDRPOINTER_REG_13__SCAN_IN & ~new_n2240_ & ~P1_STATEBS16_REG_SCAN_IN) | P1_STATE2_REG_2__SCAN_IN | (~P1_PHYADDRPOINTER_REG_13__SCAN_IN & (new_n2240_ | P1_STATEBS16_REG_SCAN_IN)));
  assign new_n2240_ = P1_PHYADDRPOINTER_REG_12__SCAN_IN & P1_PHYADDRPOINTER_REG_11__SCAN_IN & P1_PHYADDRPOINTER_REG_10__SCAN_IN & P1_PHYADDRPOINTER_REG_9__SCAN_IN & P1_PHYADDRPOINTER_REG_8__SCAN_IN & new_n2241_ & P1_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign new_n2241_ = P1_PHYADDRPOINTER_REG_6__SCAN_IN & P1_PHYADDRPOINTER_REG_5__SCAN_IN & P1_PHYADDRPOINTER_REG_4__SCAN_IN & P1_PHYADDRPOINTER_REG_3__SCAN_IN & P1_PHYADDRPOINTER_REG_2__SCAN_IN & P1_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign new_n2242_ = new_n2239_ & (~new_n2237_ | ((~new_n2227_ ^ ~new_n2163_) & new_n2047_ & (new_n2232_ ^ new_n2163_)) | ((~new_n2227_ | new_n2163_) & (new_n2227_ | ~new_n2163_) & (~new_n2047_ | (~new_n2232_ ^ new_n2163_))));
  assign new_n2243_ = ~new_n2245_ & new_n2237_ & (~new_n2047_ | new_n2244_) & (new_n2047_ | ~new_n2244_);
  assign new_n2244_ = new_n2232_ ^ ~new_n2163_;
  assign new_n2245_ = (new_n2246_ | P1_STATEBS16_REG_SCAN_IN | P1_STATE2_REG_2__SCAN_IN) & (~P1_PHYADDRPOINTER_REG_12__SCAN_IN | ~P1_STATEBS16_REG_SCAN_IN | P1_STATE2_REG_2__SCAN_IN) & (~P1_EAX_REG_12__SCAN_IN | ~new_n2053_ | ~P1_STATE2_REG_2__SCAN_IN);
  assign new_n2246_ = P1_PHYADDRPOINTER_REG_12__SCAN_IN ^ (P1_PHYADDRPOINTER_REG_11__SCAN_IN & P1_PHYADDRPOINTER_REG_10__SCAN_IN & new_n2247_ & P1_PHYADDRPOINTER_REG_9__SCAN_IN);
  assign new_n2247_ = P1_PHYADDRPOINTER_REG_8__SCAN_IN & new_n2241_ & P1_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign new_n2248_ = new_n2245_ & (~new_n2237_ | (new_n2047_ & ~new_n2244_) | (~new_n2047_ & new_n2244_));
  assign new_n2249_ = new_n2297_ & new_n2300_ & ((new_n2250_ & ~new_n2303_) | ((new_n2256_ | ~new_n2260_) & ~new_n2296_ & (new_n2250_ | ~new_n2303_)));
  assign new_n2250_ = new_n2237_ & (~new_n2252_ | (new_n2251_ & ~new_n2198_)) & ~new_n2255_ & (~new_n2253_ | (~new_n2251_ & ~new_n2185_));
  assign new_n2251_ = ~new_n2192_ & (new_n2201_ | (~new_n2049_ & (new_n2147_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_))))));
  assign new_n2252_ = new_n2177_ & (~new_n2163_ | new_n2184_);
  assign new_n2253_ = ~new_n2254_ & ~new_n2198_ & ~new_n2199_;
  assign new_n2254_ = new_n2163_ ^ ~new_n2184_;
  assign new_n2255_ = new_n2254_ ? new_n2199_ : new_n2178_;
  assign new_n2256_ = ~new_n2258_ & new_n2237_ & (~new_n2257_ | (~new_n2198_ & (new_n2251_ | new_n2185_))) & (new_n2257_ | new_n2198_ | (~new_n2251_ & ~new_n2185_));
  assign new_n2257_ = ~new_n2178_ & ~new_n2199_;
  assign new_n2258_ = (~P1_EAX_REG_6__SCAN_IN | ~new_n2053_ | ~P1_STATE2_REG_2__SCAN_IN) & (~P1_PHYADDRPOINTER_REG_6__SCAN_IN | ~P1_STATEBS16_REG_SCAN_IN | P1_STATE2_REG_2__SCAN_IN) & (new_n2259_ | P1_STATEBS16_REG_SCAN_IN | P1_STATE2_REG_2__SCAN_IN);
  assign new_n2259_ = P1_PHYADDRPOINTER_REG_6__SCAN_IN ^ (P1_PHYADDRPOINTER_REG_5__SCAN_IN & P1_PHYADDRPOINTER_REG_4__SCAN_IN & P1_PHYADDRPOINTER_REG_3__SCAN_IN & P1_PHYADDRPOINTER_REG_2__SCAN_IN & P1_PHYADDRPOINTER_REG_1__SCAN_IN);
  assign new_n2260_ = ((~new_n2263_ & (~new_n2261_ | ~new_n2237_)) | (~new_n2269_ & ~new_n2271_) | ((new_n2278_ | ~new_n2276_ | ~new_n2237_) & (~new_n2282_ | (new_n2278_ & (~new_n2276_ | ~new_n2237_))))) & (~new_n2269_ | ~new_n2271_ | (~new_n2263_ & (~new_n2261_ | ~new_n2237_))) & (~new_n2263_ | ~new_n2261_ | ~new_n2237_);
  assign new_n2261_ = ~new_n2262_ ^ (~new_n2192_ & (new_n2201_ | (~new_n2049_ & (new_n2147_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))))));
  assign new_n2262_ = ~new_n2185_ & ~new_n2198_;
  assign new_n2263_ = ((~new_n2267_ & P1_PHYADDRPOINTER_REG_5__SCAN_IN) | P1_STATE2_REG_2__SCAN_IN | (new_n2267_ & ~P1_PHYADDRPOINTER_REG_5__SCAN_IN)) & ((new_n2264_ & ~new_n2238_) | ~P1_STATE2_REG_2__SCAN_IN | (new_n2053_ & P1_EAX_REG_5__SCAN_IN));
  assign new_n2264_ = new_n2265_ & ~new_n2133_ & ~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)));
  assign new_n2265_ = new_n2266_ & new_n2137_ & P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign new_n2266_ = ~new_n2097_ & new_n2091_ & ~new_n2065_ & new_n2079_ & ~new_n2053_ & ~new_n2085_;
  assign new_n2267_ = ~P1_STATEBS16_REG_SCAN_IN & (~P1_PHYADDRPOINTER_REG_4__SCAN_IN | ~new_n2268_ | ~P1_PHYADDRPOINTER_REG_3__SCAN_IN);
  assign new_n2268_ = P1_PHYADDRPOINTER_REG_2__SCAN_IN & P1_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign new_n2269_ = new_n2237_ & (~new_n2270_ ^ (~new_n2049_ & (new_n2147_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_))))));
  assign new_n2270_ = ~new_n2201_ & ~new_n2192_;
  assign new_n2271_ = (~new_n2275_ | (new_n2272_ & (~P1_PHYADDRPOINTER_REG_4__SCAN_IN ^ (new_n2268_ & P1_PHYADDRPOINTER_REG_3__SCAN_IN)))) & (~new_n2272_ | new_n2275_ | (new_n2274_ & P1_PHYADDRPOINTER_REG_4__SCAN_IN));
  assign new_n2272_ = new_n2273_ & (~new_n2237_ | (new_n2265_ & ~new_n2133_ & ~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))) | (~new_n2265_ & (new_n2133_ | new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_))))));
  assign new_n2273_ = (~P1_EAX_REG_4__SCAN_IN | ~new_n2053_ | ~P1_STATE2_REG_2__SCAN_IN) & (~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~P1_STATE2_REG_2__SCAN_IN | new_n2053_ | new_n2085_);
  assign new_n2274_ = P1_STATEBS16_REG_SCAN_IN & ~P1_STATE2_REG_2__SCAN_IN;
  assign new_n2275_ = ~P1_STATEBS16_REG_SCAN_IN & ~P1_STATE2_REG_2__SCAN_IN;
  assign new_n2276_ = ~new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)));
  assign new_n2277_ = ~new_n2135_ ^ (new_n2145_ | (~P1_STATE2_REG_0__SCAN_IN & (new_n2133_ | new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_)))) & (~new_n2133_ | (~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))))));
  assign new_n2278_ = new_n2279_ ? ~new_n2281_ : new_n2275_;
  assign new_n2279_ = new_n2280_ & (~new_n2237_ | (~new_n2133_ & ~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))) | (new_n2133_ & (new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_))))));
  assign new_n2280_ = (~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_STATE2_REG_2__SCAN_IN | new_n2053_ | new_n2085_) & (~P1_EAX_REG_3__SCAN_IN | ~new_n2053_ | ~P1_STATE2_REG_2__SCAN_IN) & ((~new_n2268_ & ~P1_PHYADDRPOINTER_REG_3__SCAN_IN) | (new_n2268_ & P1_PHYADDRPOINTER_REG_3__SCAN_IN) | P1_STATEBS16_REG_SCAN_IN | P1_STATE2_REG_2__SCAN_IN);
  assign new_n2281_ = ~P1_STATE2_REG_2__SCAN_IN & (~P1_STATEBS16_REG_SCAN_IN | P1_PHYADDRPOINTER_REG_3__SCAN_IN);
  assign new_n2282_ = (new_n2274_ | (new_n2237_ & (~new_n2154_ | new_n2283_) & (new_n2154_ | ~new_n2283_)) | ((~new_n2285_ | (new_n2284_ & new_n2237_)) & (~new_n2287_ | (~new_n2285_ & new_n2284_ & new_n2237_)))) & (new_n2293_ | ((new_n2274_ | (new_n2237_ & (~new_n2154_ | new_n2283_) & (new_n2154_ | ~new_n2283_))) & (~new_n2285_ | (new_n2284_ & new_n2237_)) & (~new_n2287_ | (~new_n2285_ & new_n2284_ & new_n2237_))));
  assign new_n2283_ = ~new_n2200_ ^ ((~P1_STATE2_REG_0__SCAN_IN & (new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_)))) & (~new_n2131_ | (~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))) | (~new_n2149_ & new_n2079_ & P1_STATE2_REG_0__SCAN_IN));
  assign new_n2284_ = (new_n2163_ | (~new_n2156_ & ~new_n2176_) | (~new_n2175_ ^ (new_n2169_ | (~P1_STATE2_REG_0__SCAN_IN & (~new_n2121_ ^ ~new_n2155_))))) & ((~new_n2175_ & (new_n2169_ | (~P1_STATE2_REG_0__SCAN_IN & (~new_n2121_ ^ ~new_n2155_)))) | (~new_n2163_ & (new_n2156_ | new_n2176_)) | (new_n2175_ & ~new_n2169_ & (P1_STATE2_REG_0__SCAN_IN | (new_n2121_ ^ ~new_n2155_))));
  assign new_n2285_ = P1_STATE2_REG_2__SCAN_IN ? (new_n2286_ & (new_n2238_ | (new_n2121_ ^ ~new_n2155_))) : ~P1_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign new_n2286_ = (~new_n2053_ | ~P1_EAX_REG_1__SCAN_IN) & (~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | new_n2053_ | new_n2085_);
  assign new_n2287_ = (P1_PHYADDRPOINTER_REG_0__SCAN_IN | P1_STATEBS16_REG_SCAN_IN | P1_STATE2_REG_2__SCAN_IN) & (new_n2289_ | ~P1_STATE2_REG_2__SCAN_IN | ((~new_n2156_ ^ ~new_n2288_) & ~new_n2053_ & new_n2085_));
  assign new_n2288_ = ~new_n2163_ & ~new_n2176_;
  assign new_n2289_ = new_n2290_ & (new_n2238_ | (~new_n2122_ & (new_n2130_ | (P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & (new_n2127_ | ~new_n2051_ | ~new_n2128_)))) | (new_n2122_ & ~new_n2130_ & (~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~new_n2127_ & new_n2051_ & new_n2128_))));
  assign new_n2290_ = (~new_n2291_ | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~new_n2292_ | ~P1_EAX_REG_0__SCAN_IN);
  assign new_n2291_ = ~new_n2053_ & ~new_n2085_;
  assign new_n2292_ = new_n2053_ & P1_STATE2_REG_2__SCAN_IN;
  assign new_n2293_ = ~new_n2295_ & (~new_n2294_ | (~new_n2238_ & (new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_)))) & (~new_n2131_ | (~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))));
  assign new_n2294_ = (~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | new_n2053_ | new_n2085_) & P1_STATE2_REG_2__SCAN_IN & (~new_n2053_ | ~P1_EAX_REG_2__SCAN_IN);
  assign new_n2295_ = (P1_PHYADDRPOINTER_REG_2__SCAN_IN | P1_STATEBS16_REG_SCAN_IN | P1_PHYADDRPOINTER_REG_1__SCAN_IN) & ~P1_STATE2_REG_2__SCAN_IN & (~P1_PHYADDRPOINTER_REG_2__SCAN_IN | (~P1_STATEBS16_REG_SCAN_IN & ~P1_PHYADDRPOINTER_REG_1__SCAN_IN));
  assign new_n2296_ = new_n2258_ & (~new_n2237_ | (new_n2257_ & (new_n2198_ | (~new_n2251_ & ~new_n2185_))) | (~new_n2257_ & ~new_n2198_ & (new_n2251_ | new_n2185_)));
  assign new_n2297_ = (~new_n2298_ | (new_n2237_ & (new_n2202_ | new_n2209_ | new_n2215_ | new_n2048_ | new_n2221_) & (~new_n2202_ | (~new_n2209_ & ~new_n2215_ & ~new_n2048_ & ~new_n2221_)))) & (~new_n2299_ | (new_n2237_ & (new_n2209_ | new_n2215_ | new_n2048_ | new_n2221_) & (~new_n2209_ | (~new_n2215_ & ~new_n2048_ & ~new_n2221_))));
  assign new_n2298_ = (~P1_EAX_REG_11__SCAN_IN | ~new_n2053_ | ~P1_STATE2_REG_2__SCAN_IN) & ((P1_PHYADDRPOINTER_REG_11__SCAN_IN & ~P1_STATEBS16_REG_SCAN_IN & (~P1_PHYADDRPOINTER_REG_10__SCAN_IN | ~new_n2247_ | ~P1_PHYADDRPOINTER_REG_9__SCAN_IN)) | P1_STATE2_REG_2__SCAN_IN | (~P1_PHYADDRPOINTER_REG_11__SCAN_IN & (P1_STATEBS16_REG_SCAN_IN | (P1_PHYADDRPOINTER_REG_10__SCAN_IN & new_n2247_ & P1_PHYADDRPOINTER_REG_9__SCAN_IN))));
  assign new_n2299_ = (~P1_EAX_REG_10__SCAN_IN | ~new_n2053_ | ~P1_STATE2_REG_2__SCAN_IN) & ((P1_PHYADDRPOINTER_REG_10__SCAN_IN & ~P1_STATEBS16_REG_SCAN_IN & (~new_n2247_ | ~P1_PHYADDRPOINTER_REG_9__SCAN_IN)) | P1_STATE2_REG_2__SCAN_IN | (~P1_PHYADDRPOINTER_REG_10__SCAN_IN & (P1_STATEBS16_REG_SCAN_IN | (new_n2247_ & P1_PHYADDRPOINTER_REG_9__SCAN_IN))));
  assign new_n2300_ = (~new_n2301_ | (new_n2237_ & (new_n2215_ | new_n2048_ | new_n2221_) & (~new_n2215_ | (~new_n2048_ & ~new_n2221_)))) & (~new_n2302_ | (new_n2237_ & (~new_n2048_ | ~new_n2221_) & (new_n2048_ | new_n2221_)));
  assign new_n2301_ = (~P1_EAX_REG_9__SCAN_IN | ~new_n2053_ | ~P1_STATE2_REG_2__SCAN_IN) & ((P1_PHYADDRPOINTER_REG_9__SCAN_IN & ~new_n2247_ & ~P1_STATEBS16_REG_SCAN_IN) | P1_STATE2_REG_2__SCAN_IN | (~P1_PHYADDRPOINTER_REG_9__SCAN_IN & (new_n2247_ | P1_STATEBS16_REG_SCAN_IN)));
  assign new_n2302_ = (~P1_EAX_REG_8__SCAN_IN | ~new_n2053_ | ~P1_STATE2_REG_2__SCAN_IN) & ((P1_PHYADDRPOINTER_REG_8__SCAN_IN & ~P1_STATEBS16_REG_SCAN_IN & (~new_n2241_ | ~P1_PHYADDRPOINTER_REG_7__SCAN_IN)) | P1_STATE2_REG_2__SCAN_IN | (~P1_PHYADDRPOINTER_REG_8__SCAN_IN & (P1_STATEBS16_REG_SCAN_IN | (new_n2241_ & P1_PHYADDRPOINTER_REG_7__SCAN_IN))));
  assign new_n2303_ = (~P1_EAX_REG_7__SCAN_IN | ~new_n2053_ | ~P1_STATE2_REG_2__SCAN_IN) & ((P1_PHYADDRPOINTER_REG_7__SCAN_IN & ~new_n2241_ & ~P1_STATEBS16_REG_SCAN_IN) | P1_STATE2_REG_2__SCAN_IN | (~P1_PHYADDRPOINTER_REG_7__SCAN_IN & (new_n2241_ | P1_STATEBS16_REG_SCAN_IN)));
  assign new_n2304_ = (new_n2298_ | ~new_n2237_ | (new_n2305_ & (~new_n2203_ ^ ~new_n2163_)) | (~new_n2305_ & (~new_n2203_ | new_n2163_) & (new_n2203_ | ~new_n2163_))) & ((new_n2298_ & (~new_n2237_ | (new_n2305_ & (~new_n2203_ ^ ~new_n2163_)) | (~new_n2305_ & (~new_n2203_ | new_n2163_) & (new_n2203_ | ~new_n2163_)))) | (new_n2299_ & (~new_n2306_ | ~new_n2237_)) | (new_n2307_ & (new_n2299_ | ~new_n2306_ | ~new_n2237_)));
  assign new_n2305_ = ~new_n2209_ & ~new_n2215_ & ~new_n2048_ & ~new_n2221_;
  assign new_n2306_ = ~new_n2209_ ^ (~new_n2215_ & ~new_n2048_ & ~new_n2221_);
  assign new_n2307_ = ((new_n2301_ & (~new_n2237_ | (~new_n2215_ & ~new_n2048_ & ~new_n2221_) | (new_n2215_ & (new_n2048_ | new_n2221_)))) | new_n2302_ | ~new_n2237_ | (new_n2048_ & new_n2221_) | (~new_n2048_ & ~new_n2221_)) & (new_n2301_ | ~new_n2237_ | (~new_n2215_ & ~new_n2048_ & ~new_n2221_) | (new_n2215_ & (new_n2048_ | new_n2221_)));
  assign new_n2308_ = (~new_n2321_ | (new_n2237_ & ((~new_n2316_ ^ new_n2163_) | ~new_n2309_ | (new_n2311_ ^ ~new_n2163_)) & ((~new_n2316_ & new_n2163_) | (new_n2316_ & ~new_n2163_) | (new_n2309_ & (~new_n2311_ ^ ~new_n2163_))))) & (~new_n2322_ | (new_n2237_ & (~new_n2309_ | (new_n2311_ ^ ~new_n2163_)) & (new_n2309_ | (new_n2311_ & ~new_n2163_) | (~new_n2311_ & new_n2163_))));
  assign new_n2309_ = ~new_n2310_ & ~new_n2244_ & ~new_n2202_ & ~new_n2209_ & ~new_n2215_ & ~new_n2048_ & ~new_n2221_;
  assign new_n2310_ = new_n2227_ ^ ~new_n2163_;
  assign new_n2311_ = ~new_n2204_ & (~new_n2312_ | ~new_n2313_ | ~new_n2315_ | (new_n2056_ & P1_INSTQUEUE_REG_1__6__SCAN_IN) | (new_n2080_ & P1_INSTQUEUE_REG_9__6__SCAN_IN));
  assign new_n2312_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_5__6__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_13__6__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_8__6__SCAN_IN);
  assign new_n2313_ = new_n2314_ & (~P1_INSTQUEUE_REG_15__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_6__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2314_ = (~P1_INSTQUEUE_REG_4__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_0__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2315_ = (~P1_INSTQUEUE_REG_2__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_14__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2316_ = ~new_n2204_ & (~new_n2317_ | ~new_n2318_ | ~new_n2320_ | (new_n2056_ & P1_INSTQUEUE_REG_1__7__SCAN_IN) | (new_n2080_ & P1_INSTQUEUE_REG_9__7__SCAN_IN));
  assign new_n2317_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_5__7__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_13__7__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_8__7__SCAN_IN);
  assign new_n2318_ = new_n2319_ & (~P1_INSTQUEUE_REG_15__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_6__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2319_ = (~P1_INSTQUEUE_REG_4__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_0__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2320_ = (~P1_INSTQUEUE_REG_2__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_14__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_10__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2321_ = (~P1_EAX_REG_15__SCAN_IN | ~new_n2053_ | ~P1_STATE2_REG_2__SCAN_IN) & ((P1_PHYADDRPOINTER_REG_15__SCAN_IN & ~P1_STATEBS16_REG_SCAN_IN & (~P1_PHYADDRPOINTER_REG_14__SCAN_IN | ~new_n2240_ | ~P1_PHYADDRPOINTER_REG_13__SCAN_IN)) | P1_STATE2_REG_2__SCAN_IN | (~P1_PHYADDRPOINTER_REG_15__SCAN_IN & (P1_STATEBS16_REG_SCAN_IN | (P1_PHYADDRPOINTER_REG_14__SCAN_IN & new_n2240_ & P1_PHYADDRPOINTER_REG_13__SCAN_IN))));
  assign new_n2322_ = (P1_STATEBS16_REG_SCAN_IN | P1_STATE2_REG_2__SCAN_IN | (P1_PHYADDRPOINTER_REG_14__SCAN_IN ^ (new_n2240_ & P1_PHYADDRPOINTER_REG_13__SCAN_IN))) & (~P1_EAX_REG_14__SCAN_IN | ~new_n2053_ | ~P1_STATE2_REG_2__SCAN_IN) & (~P1_PHYADDRPOINTER_REG_14__SCAN_IN | ~P1_STATEBS16_REG_SCAN_IN | P1_STATE2_REG_2__SCAN_IN);
  assign new_n2323_ = (new_n2321_ | ~new_n2237_ | ((new_n2316_ ^ new_n2163_) & new_n2309_ & (~new_n2311_ ^ ~new_n2163_)) | ((new_n2316_ | ~new_n2163_) & (~new_n2316_ | new_n2163_) & (~new_n2309_ | (new_n2311_ ^ ~new_n2163_)))) & ((new_n2321_ & (~new_n2237_ | ((new_n2316_ ^ new_n2163_) & new_n2309_ & (~new_n2311_ ^ ~new_n2163_)) | ((new_n2316_ | ~new_n2163_) & (~new_n2316_ | new_n2163_) & (~new_n2309_ | (new_n2311_ ^ ~new_n2163_))))) | new_n2322_ | ~new_n2237_ | (new_n2309_ & (~new_n2311_ ^ ~new_n2163_)) | (~new_n2309_ & (~new_n2311_ | new_n2163_) & (new_n2311_ | ~new_n2163_)));
  assign new_n2324_ = new_n2237_ & new_n2163_ & (~new_n2325_ | (~new_n2316_ ^ new_n2163_));
  assign new_n2325_ = ~new_n2326_ & ~new_n2310_ & ~new_n2244_ & ~new_n2202_ & ~new_n2209_ & ~new_n2215_ & ~new_n2048_ & ~new_n2221_;
  assign new_n2326_ = new_n2311_ ^ ~new_n2163_;
  assign new_n2327_ = new_n2328_ & new_n2237_ & ((new_n2163_ & (~new_n2325_ | (~new_n2316_ ^ new_n2163_))) | (new_n2325_ & new_n2316_ & ~new_n2163_));
  assign new_n2328_ = new_n2329_ ? (new_n2275_ & (~P1_PHYADDRPOINTER_REG_16__SCAN_IN ^ (P1_PHYADDRPOINTER_REG_15__SCAN_IN & P1_PHYADDRPOINTER_REG_14__SCAN_IN & new_n2240_ & P1_PHYADDRPOINTER_REG_13__SCAN_IN))) : ~new_n2275_;
  assign new_n2329_ = (~new_n2330_ | new_n2333_) & (~new_n2274_ | ~P1_PHYADDRPOINTER_REG_16__SCAN_IN) & (~new_n2292_ | ~P1_EAX_REG_16__SCAN_IN);
  assign new_n2330_ = new_n2237_ & new_n2331_;
  assign new_n2331_ = ~new_n2332_ & P1_STATE2_REG_0__SCAN_IN;
  assign new_n2332_ = (~new_n2067_ | ~new_n2073_ | ~new_n2097_ | new_n2065_ | new_n2053_ | new_n2079_ | ~new_n2085_) & (new_n2073_ | new_n2091_ | new_n2067_ | ~new_n2097_ | new_n2065_ | new_n2053_ | new_n2079_ | ~new_n2085_);
  assign new_n2333_ = new_n2334_ & new_n2335_ & new_n2337_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_2__0__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_9__0__SCAN_IN);
  assign new_n2334_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_6__0__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_14__0__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_10__0__SCAN_IN);
  assign new_n2335_ = new_n2336_ & (~P1_INSTQUEUE_REG_12__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_13__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_8__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2336_ = (~P1_INSTQUEUE_REG_11__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_1__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_0__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_4__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2337_ = (~P1_INSTQUEUE_REG_5__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_15__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2338_ = ~new_n2328_ & (~new_n2237_ | ((~new_n2163_ | (new_n2325_ & (new_n2316_ ^ new_n2163_))) & (~new_n2325_ | ~new_n2316_ | new_n2163_)));
  assign new_n2339_ = new_n2340_ ? (~new_n2275_ | (P1_PHYADDRPOINTER_REG_17__SCAN_IN ^ (P1_PHYADDRPOINTER_REG_16__SCAN_IN & P1_PHYADDRPOINTER_REG_15__SCAN_IN & P1_PHYADDRPOINTER_REG_14__SCAN_IN & new_n2240_ & P1_PHYADDRPOINTER_REG_13__SCAN_IN))) : new_n2275_;
  assign new_n2340_ = (~new_n2330_ | new_n2341_) & (~new_n2274_ | ~P1_PHYADDRPOINTER_REG_17__SCAN_IN) & (~new_n2292_ | ~P1_EAX_REG_17__SCAN_IN);
  assign new_n2341_ = new_n2342_ & new_n2343_ & new_n2345_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_2__1__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_9__1__SCAN_IN);
  assign new_n2342_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_6__1__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_14__1__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_10__1__SCAN_IN);
  assign new_n2343_ = new_n2344_ & (~P1_INSTQUEUE_REG_12__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_13__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_8__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2344_ = (~P1_INSTQUEUE_REG_0__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_4__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_1__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2345_ = (~P1_INSTQUEUE_REG_5__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_15__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2346_ = ((~new_n2330_ | new_n2348_) & (~P1_EAX_REG_18__SCAN_IN | ~new_n2053_ | ~P1_STATE2_REG_2__SCAN_IN) & (~P1_PHYADDRPOINTER_REG_18__SCAN_IN | ~P1_STATEBS16_REG_SCAN_IN | P1_STATE2_REG_2__SCAN_IN)) ? ((new_n2347_ ^ ~P1_PHYADDRPOINTER_REG_18__SCAN_IN) & ~P1_STATEBS16_REG_SCAN_IN & ~P1_STATE2_REG_2__SCAN_IN) : (P1_STATEBS16_REG_SCAN_IN | P1_STATE2_REG_2__SCAN_IN);
  assign new_n2347_ = P1_PHYADDRPOINTER_REG_17__SCAN_IN & P1_PHYADDRPOINTER_REG_16__SCAN_IN & P1_PHYADDRPOINTER_REG_15__SCAN_IN & P1_PHYADDRPOINTER_REG_14__SCAN_IN & new_n2240_ & P1_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign new_n2348_ = new_n2349_ & new_n2350_ & new_n2352_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_2__2__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_9__2__SCAN_IN);
  assign new_n2349_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_6__2__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_14__2__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_10__2__SCAN_IN);
  assign new_n2350_ = new_n2351_ & (~P1_INSTQUEUE_REG_12__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_13__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_8__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2351_ = (~P1_INSTQUEUE_REG_0__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_4__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_1__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2352_ = (~P1_INSTQUEUE_REG_5__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_15__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2353_ = ((~P1_STATEBS16_REG_SCAN_IN & ~P1_STATE2_REG_2__SCAN_IN) | ((~new_n2330_ | new_n2355_) & (~P1_EAX_REG_20__SCAN_IN | ~new_n2053_ | ~P1_STATE2_REG_2__SCAN_IN) & (~P1_PHYADDRPOINTER_REG_20__SCAN_IN | ~P1_STATEBS16_REG_SCAN_IN | P1_STATE2_REG_2__SCAN_IN))) & ((~new_n2354_ ^ ~P1_PHYADDRPOINTER_REG_20__SCAN_IN) | P1_STATEBS16_REG_SCAN_IN | P1_STATE2_REG_2__SCAN_IN | (new_n2330_ & ~new_n2355_) | (P1_EAX_REG_20__SCAN_IN & new_n2053_ & P1_STATE2_REG_2__SCAN_IN) | (P1_PHYADDRPOINTER_REG_20__SCAN_IN & P1_STATEBS16_REG_SCAN_IN & ~P1_STATE2_REG_2__SCAN_IN));
  assign new_n2354_ = P1_PHYADDRPOINTER_REG_19__SCAN_IN & P1_PHYADDRPOINTER_REG_18__SCAN_IN & P1_PHYADDRPOINTER_REG_17__SCAN_IN & P1_PHYADDRPOINTER_REG_16__SCAN_IN & P1_PHYADDRPOINTER_REG_15__SCAN_IN & P1_PHYADDRPOINTER_REG_14__SCAN_IN & new_n2240_ & P1_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign new_n2355_ = new_n2356_ & new_n2357_ & new_n2359_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_2__4__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_9__4__SCAN_IN);
  assign new_n2356_ = (~new_n2057_ | ~P1_INSTQUEUE_REG_14__4__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_10__4__SCAN_IN) & (~new_n2099_ | ~P1_INSTQUEUE_REG_6__4__SCAN_IN);
  assign new_n2357_ = new_n2358_ & (~P1_INSTQUEUE_REG_12__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_7__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_8__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2358_ = (~P1_INSTQUEUE_REG_1__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_0__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_13__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2359_ = (~P1_INSTQUEUE_REG_3__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_4__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_15__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_5__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2360_ = ((~new_n2330_ | new_n2361_) & (~new_n2274_ | ~P1_PHYADDRPOINTER_REG_19__SCAN_IN) & (~new_n2292_ | ~P1_EAX_REG_19__SCAN_IN)) ? (~new_n2366_ & new_n2275_) : ~new_n2275_;
  assign new_n2361_ = new_n2362_ & new_n2363_ & new_n2365_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_2__3__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_9__3__SCAN_IN);
  assign new_n2362_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_6__3__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_14__3__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_10__3__SCAN_IN);
  assign new_n2363_ = new_n2364_ & (~P1_INSTQUEUE_REG_12__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_13__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_8__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2364_ = (~P1_INSTQUEUE_REG_0__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_4__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_1__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2365_ = (~P1_INSTQUEUE_REG_5__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_15__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2366_ = P1_PHYADDRPOINTER_REG_19__SCAN_IN ^ (P1_PHYADDRPOINTER_REG_18__SCAN_IN & P1_PHYADDRPOINTER_REG_17__SCAN_IN & P1_PHYADDRPOINTER_REG_16__SCAN_IN & P1_PHYADDRPOINTER_REG_15__SCAN_IN & P1_PHYADDRPOINTER_REG_14__SCAN_IN & new_n2240_ & P1_PHYADDRPOINTER_REG_13__SCAN_IN);
  assign new_n2367_ = (~new_n2324_ | new_n2390_) & new_n2368_ & (~new_n2324_ | new_n2419_);
  assign new_n2368_ = (~new_n2324_ | ~new_n2369_) & (~new_n2324_ | new_n2382_);
  assign new_n2369_ = (~new_n2370_ & (~new_n2274_ | ~P1_PHYADDRPOINTER_REG_23__SCAN_IN) & (~new_n2292_ | ~P1_EAX_REG_23__SCAN_IN)) ? (new_n2275_ & (new_n2381_ ^ ~P1_PHYADDRPOINTER_REG_23__SCAN_IN)) : ~new_n2275_;
  assign new_n2370_ = (~new_n2331_ | new_n2371_ | new_n2376_) & (~new_n2371_ | ~new_n2376_) & new_n2237_ & new_n2331_;
  assign new_n2371_ = new_n2372_ & new_n2373_ & new_n2375_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_3__0__SCAN_IN) & (~new_n2099_ | ~P1_INSTQUEUE_REG_7__0__SCAN_IN);
  assign new_n2372_ = (~new_n2098_ | ~P1_INSTQUEUE_REG_10__0__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_15__0__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_11__0__SCAN_IN);
  assign new_n2373_ = new_n2374_ & (~P1_INSTQUEUE_REG_0__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_1__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2374_ = (~P1_INSTQUEUE_REG_13__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_2__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_4__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2375_ = (~P1_INSTQUEUE_REG_9__0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_6__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_8__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_5__0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2376_ = new_n2377_ & new_n2378_ & new_n2380_ & (~new_n2080_ | ~P1_INSTQUEUE_REG_10__7__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_9__7__SCAN_IN);
  assign new_n2377_ = (~new_n2099_ | ~P1_INSTQUEUE_REG_6__7__SCAN_IN) & (~new_n2056_ | ~P1_INSTQUEUE_REG_2__7__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_14__7__SCAN_IN);
  assign new_n2378_ = new_n2379_ & (~P1_INSTQUEUE_REG_13__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_1__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_15__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2379_ = (~P1_INSTQUEUE_REG_12__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_7__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_0__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2380_ = (~P1_INSTQUEUE_REG_4__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_11__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_5__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_8__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2381_ = P1_PHYADDRPOINTER_REG_22__SCAN_IN & P1_PHYADDRPOINTER_REG_21__SCAN_IN & new_n2354_ & P1_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign new_n2382_ = (new_n2383_ | new_n2275_) & (~new_n2383_ | ~new_n2275_ | (P1_PHYADDRPOINTER_REG_24__SCAN_IN ^ (new_n2381_ & P1_PHYADDRPOINTER_REG_23__SCAN_IN)));
  assign new_n2383_ = (((~new_n2331_ | new_n2385_) & (~new_n2331_ | ~new_n2384_)) | ~new_n2237_ | (~new_n2385_ & new_n2331_ & new_n2384_)) & (~new_n2292_ | ~P1_EAX_REG_24__SCAN_IN) & (~new_n2274_ | ~P1_PHYADDRPOINTER_REG_24__SCAN_IN);
  assign new_n2384_ = ~new_n2371_ & ~new_n2376_;
  assign new_n2385_ = new_n2386_ & new_n2387_ & new_n2389_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_3__1__SCAN_IN) & (~new_n2099_ | ~P1_INSTQUEUE_REG_7__1__SCAN_IN);
  assign new_n2386_ = (~new_n2098_ | ~P1_INSTQUEUE_REG_10__1__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_15__1__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_11__1__SCAN_IN);
  assign new_n2387_ = new_n2388_ & (~P1_INSTQUEUE_REG_0__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_1__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2388_ = (~P1_INSTQUEUE_REG_2__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_12__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_4__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2389_ = (~P1_INSTQUEUE_REG_9__1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_6__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_8__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_5__1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2390_ = (new_n2391_ | new_n2275_) & (~new_n2391_ | ~new_n2275_ | (P1_PHYADDRPOINTER_REG_28__SCAN_IN ^ (new_n2418_ & P1_PHYADDRPOINTER_REG_27__SCAN_IN))) & new_n2414_ & (new_n2417_ | new_n2275_) & (~new_n2417_ | ~new_n2275_ | (new_n2418_ ^ P1_PHYADDRPOINTER_REG_27__SCAN_IN));
  assign new_n2391_ = (~new_n2292_ | ~P1_EAX_REG_28__SCAN_IN) & (~new_n2274_ | ~P1_PHYADDRPOINTER_REG_28__SCAN_IN) & ((~new_n2392_ & (~new_n2331_ | new_n2409_)) | ~new_n2237_ | (new_n2392_ & ~new_n2409_));
  assign new_n2392_ = new_n2393_ & new_n2404_;
  assign new_n2393_ = ~new_n2399_ & new_n2331_ & ~new_n2394_ & ~new_n2385_ & new_n2384_;
  assign new_n2394_ = new_n2395_ & new_n2396_ & new_n2398_ & (~new_n2057_ | ~P1_INSTQUEUE_REG_15__2__SCAN_IN) & (~new_n2099_ | ~P1_INSTQUEUE_REG_7__2__SCAN_IN);
  assign new_n2395_ = (~new_n2098_ | ~P1_INSTQUEUE_REG_10__2__SCAN_IN) & (~new_n2056_ | ~P1_INSTQUEUE_REG_3__2__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_11__2__SCAN_IN);
  assign new_n2396_ = new_n2397_ & (~P1_INSTQUEUE_REG_4__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_0__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_12__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2397_ = (~P1_INSTQUEUE_REG_8__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_6__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_2__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2398_ = (~P1_INSTQUEUE_REG_9__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_5__2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_1__2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2399_ = new_n2400_ & new_n2401_ & new_n2403_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_3__3__SCAN_IN) & (~new_n2099_ | ~P1_INSTQUEUE_REG_7__3__SCAN_IN);
  assign new_n2400_ = (~new_n2098_ | ~P1_INSTQUEUE_REG_10__3__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_15__3__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_11__3__SCAN_IN);
  assign new_n2401_ = new_n2402_ & (~P1_INSTQUEUE_REG_0__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_1__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2402_ = (~P1_INSTQUEUE_REG_2__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_12__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_4__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2403_ = (~P1_INSTQUEUE_REG_9__3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_6__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_8__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_5__3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2404_ = new_n2331_ & (~new_n2405_ | ~new_n2406_ | ~new_n2408_ | (new_n2056_ & P1_INSTQUEUE_REG_3__4__SCAN_IN) | (new_n2099_ & P1_INSTQUEUE_REG_7__4__SCAN_IN));
  assign new_n2405_ = (~new_n2098_ | ~P1_INSTQUEUE_REG_10__4__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_15__4__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_11__4__SCAN_IN);
  assign new_n2406_ = new_n2407_ & (~P1_INSTQUEUE_REG_6__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_12__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2407_ = (~P1_INSTQUEUE_REG_14__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_1__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_2__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_4__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2408_ = (~P1_INSTQUEUE_REG_5__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_9__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_8__4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_0__4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2409_ = new_n2410_ & new_n2411_ & new_n2413_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_3__5__SCAN_IN) & (~new_n2099_ | ~P1_INSTQUEUE_REG_7__5__SCAN_IN);
  assign new_n2410_ = (~new_n2098_ | ~P1_INSTQUEUE_REG_10__5__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_15__5__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_11__5__SCAN_IN);
  assign new_n2411_ = new_n2412_ & (~P1_INSTQUEUE_REG_0__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_1__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2412_ = (~P1_INSTQUEUE_REG_2__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_12__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_4__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2413_ = (~P1_INSTQUEUE_REG_9__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_6__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_8__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_5__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2414_ = (new_n2415_ | new_n2275_) & (~new_n2415_ | ~new_n2275_ | (P1_PHYADDRPOINTER_REG_26__SCAN_IN ^ (P1_PHYADDRPOINTER_REG_25__SCAN_IN & P1_PHYADDRPOINTER_REG_24__SCAN_IN & new_n2381_ & P1_PHYADDRPOINTER_REG_23__SCAN_IN)));
  assign new_n2415_ = ~new_n2416_ & (~new_n2292_ | ~P1_EAX_REG_26__SCAN_IN) & (~new_n2274_ | ~P1_PHYADDRPOINTER_REG_26__SCAN_IN);
  assign new_n2416_ = ((new_n2331_ & ~new_n2399_) | (new_n2331_ & ~new_n2394_ & ~new_n2385_ & new_n2384_)) & new_n2237_ & (new_n2399_ | ~new_n2331_ | new_n2394_ | new_n2385_ | ~new_n2384_);
  assign new_n2417_ = ((~new_n2393_ & ~new_n2404_) | ~new_n2237_ | (new_n2393_ & new_n2404_)) & (~new_n2274_ | ~P1_PHYADDRPOINTER_REG_27__SCAN_IN) & (~new_n2292_ | ~P1_EAX_REG_27__SCAN_IN);
  assign new_n2418_ = P1_PHYADDRPOINTER_REG_26__SCAN_IN & P1_PHYADDRPOINTER_REG_25__SCAN_IN & P1_PHYADDRPOINTER_REG_24__SCAN_IN & P1_PHYADDRPOINTER_REG_23__SCAN_IN & P1_PHYADDRPOINTER_REG_22__SCAN_IN & P1_PHYADDRPOINTER_REG_21__SCAN_IN & new_n2354_ & P1_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign new_n2419_ = (new_n2420_ | new_n2275_) & (~new_n2420_ | ~new_n2275_ | (P1_PHYADDRPOINTER_REG_25__SCAN_IN ^ (P1_PHYADDRPOINTER_REG_24__SCAN_IN & new_n2381_ & P1_PHYADDRPOINTER_REG_23__SCAN_IN)));
  assign new_n2420_ = ~new_n2421_ & (~new_n2292_ | ~P1_EAX_REG_25__SCAN_IN) & (~new_n2274_ | ~P1_PHYADDRPOINTER_REG_25__SCAN_IN);
  assign new_n2421_ = ((new_n2331_ & ~new_n2394_) | (~new_n2385_ & new_n2331_ & new_n2384_)) & new_n2237_ & (~new_n2331_ | new_n2394_ | new_n2385_ | ~new_n2384_);
  assign new_n2422_ = (~new_n2324_ | ~new_n2360_) & (~new_n2324_ | new_n2353_);
  assign new_n2423_ = (new_n2324_ | ~new_n2382_) & (new_n2324_ | new_n2369_);
  assign new_n2424_ = ~new_n2419_ & ~new_n2414_ & ((~new_n2417_ & ~new_n2275_) | ((new_n2418_ ^ ~P1_PHYADDRPOINTER_REG_27__SCAN_IN) & new_n2417_ & new_n2275_));
  assign new_n2425_ = new_n2426_ ? (new_n2275_ & (~P1_PHYADDRPOINTER_REG_22__SCAN_IN ^ (P1_PHYADDRPOINTER_REG_21__SCAN_IN & new_n2354_ & P1_PHYADDRPOINTER_REG_20__SCAN_IN))) : ~new_n2275_;
  assign new_n2426_ = (~new_n2330_ | new_n2427_) & (~new_n2274_ | ~P1_PHYADDRPOINTER_REG_22__SCAN_IN) & (~new_n2292_ | ~P1_EAX_REG_22__SCAN_IN);
  assign new_n2427_ = new_n2428_ & new_n2429_ & new_n2431_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_2__6__SCAN_IN) & (~new_n2098_ | ~P1_INSTQUEUE_REG_9__6__SCAN_IN);
  assign new_n2428_ = (~new_n2057_ | ~P1_INSTQUEUE_REG_14__6__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_10__6__SCAN_IN) & (~new_n2099_ | ~P1_INSTQUEUE_REG_6__6__SCAN_IN);
  assign new_n2429_ = new_n2430_ & (~P1_INSTQUEUE_REG_1__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_15__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_4__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2430_ = (~P1_INSTQUEUE_REG_8__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_13__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_5__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2431_ = (~P1_INSTQUEUE_REG_0__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_11__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2432_ = (~new_n2433_ & (~new_n2274_ | ~P1_PHYADDRPOINTER_REG_21__SCAN_IN) & (~new_n2292_ | ~P1_EAX_REG_21__SCAN_IN)) ? (~new_n2438_ & new_n2275_) : ~new_n2275_;
  assign new_n2433_ = new_n2330_ & (~new_n2434_ | ~new_n2435_ | ~new_n2437_ | (new_n2056_ & P1_INSTQUEUE_REG_2__5__SCAN_IN) | (new_n2098_ & P1_INSTQUEUE_REG_9__5__SCAN_IN));
  assign new_n2434_ = (~new_n2057_ | ~P1_INSTQUEUE_REG_14__5__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_10__5__SCAN_IN) & (~new_n2099_ | ~P1_INSTQUEUE_REG_6__5__SCAN_IN);
  assign new_n2435_ = new_n2436_ & (~P1_INSTQUEUE_REG_1__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_15__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_4__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2436_ = (~P1_INSTQUEUE_REG_8__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_13__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_5__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_12__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2437_ = (~P1_INSTQUEUE_REG_0__5__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_3__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_7__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_11__5__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2438_ = P1_PHYADDRPOINTER_REG_21__SCAN_IN ^ (new_n2354_ & P1_PHYADDRPOINTER_REG_20__SCAN_IN);
  assign new_n2439_ = new_n2324_ ^ new_n2440_;
  assign new_n2440_ = new_n2441_ ? (~new_n2448_ & new_n2275_) : ~new_n2275_;
  assign new_n2441_ = ((~new_n2442_ & ~new_n2443_) | ~new_n2237_ | (new_n2442_ & new_n2443_)) & (~new_n2274_ | ~P1_PHYADDRPOINTER_REG_29__SCAN_IN) & (~new_n2292_ | ~P1_EAX_REG_29__SCAN_IN);
  assign new_n2442_ = new_n2392_ & ~new_n2409_;
  assign new_n2443_ = new_n2331_ & (~new_n2444_ | ~new_n2445_ | ~new_n2447_ | (new_n2057_ & P1_INSTQUEUE_REG_15__6__SCAN_IN) | (new_n2099_ & P1_INSTQUEUE_REG_7__6__SCAN_IN));
  assign new_n2444_ = (~new_n2098_ | ~P1_INSTQUEUE_REG_10__6__SCAN_IN) & (~new_n2056_ | ~P1_INSTQUEUE_REG_3__6__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_11__6__SCAN_IN);
  assign new_n2445_ = new_n2446_ & (~P1_INSTQUEUE_REG_4__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_0__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_12__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2446_ = (~P1_INSTQUEUE_REG_8__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_6__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_2__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2447_ = (~P1_INSTQUEUE_REG_9__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_5__6__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_1__6__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2448_ = P1_PHYADDRPOINTER_REG_29__SCAN_IN ^ (P1_PHYADDRPOINTER_REG_28__SCAN_IN & new_n2418_ & P1_PHYADDRPOINTER_REG_27__SCAN_IN);
  assign new_n2449_ = ~new_n2324_ & (new_n2391_ | new_n2275_) & (~new_n2391_ | ~new_n2275_ | (P1_PHYADDRPOINTER_REG_28__SCAN_IN ^ (new_n2418_ & P1_PHYADDRPOINTER_REG_27__SCAN_IN)));
  assign new_n2450_ = new_n2451_ & (new_n2090_ | (new_n2456_ & P1_INSTADDRPOINTER_REG_25__SCAN_IN) | (~new_n2455_ & P1_EBX_REG_25__SCAN_IN)) & (~new_n2090_ | ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_25__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_25__SCAN_IN)));
  assign new_n2451_ = new_n2452_ & (new_n2090_ | (new_n2456_ & P1_INSTADDRPOINTER_REG_24__SCAN_IN) | (~new_n2455_ & P1_EBX_REG_24__SCAN_IN)) & (~new_n2090_ | ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_24__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_24__SCAN_IN)));
  assign new_n2452_ = new_n2475_ & new_n2472_ & ~new_n2474_ & new_n2453_ & new_n2473_;
  assign new_n2453_ = new_n2471_ & new_n2470_ & new_n2454_ & ~new_n2469_ & new_n2468_ & new_n2467_ & new_n2457_ & new_n2463_;
  assign new_n2454_ = ~new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_16__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_16__SCAN_IN));
  assign new_n2455_ = new_n2091_ ? new_n2073_ : new_n2067_;
  assign new_n2456_ = (new_n2073_ | ~new_n2116_) & (new_n2067_ | new_n2073_);
  assign new_n2457_ = ~new_n2462_ & ~new_n2461_ & ~new_n2458_ & ~new_n2459_ & ~new_n2460_;
  assign new_n2458_ = ((~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_) | ((new_n2067_ | new_n2091_) & (~P1_EBX_REG_1__SCAN_IN | (new_n2091_ ? new_n2073_ : new_n2067_)) & (~P1_INSTADDRPOINTER_REG_1__SCAN_IN | (~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_))) | (~new_n2067_ & ~new_n2091_ & ((P1_EBX_REG_1__SCAN_IN & (new_n2091_ ? ~new_n2073_ : ~new_n2067_)) | (P1_INSTADDRPOINTER_REG_1__SCAN_IN & (new_n2067_ | new_n2073_) & (new_n2073_ | ~new_n2116_))))) & (new_n2073_ | ~new_n2091_ | (~P1_EBX_REG_0__SCAN_IN & (~P1_INSTADDRPOINTER_REG_0__SCAN_IN | (~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_)))) & (new_n2067_ | new_n2091_ | P1_EBX_REG_0__SCAN_IN | (P1_INSTADDRPOINTER_REG_0__SCAN_IN & (new_n2067_ | new_n2073_) & (new_n2073_ | ~new_n2116_)));
  assign new_n2459_ = ((~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_)) & ((~new_n2067_ & ~new_n2091_) ^ ((~P1_EBX_REG_1__SCAN_IN | (new_n2091_ ? new_n2073_ : new_n2067_)) & (~P1_INSTADDRPOINTER_REG_1__SCAN_IN | (~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_))));
  assign new_n2460_ = ((~P1_INSTADDRPOINTER_REG_2__SCAN_IN | (~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_)) & (~P1_EBX_REG_2__SCAN_IN | (new_n2091_ ? new_n2073_ : new_n2067_))) ? (new_n2067_ | new_n2091_ | (P1_EBX_REG_3__SCAN_IN & (new_n2091_ ? ~new_n2073_ : ~new_n2067_)) | (P1_INSTADDRPOINTER_REG_3__SCAN_IN & (new_n2067_ | new_n2073_) & (new_n2073_ | ~new_n2116_))) : ((~new_n2067_ & ~new_n2091_) | ((~P1_EBX_REG_3__SCAN_IN | (new_n2091_ ? new_n2073_ : new_n2067_)) & (~P1_INSTADDRPOINTER_REG_3__SCAN_IN | (~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_))));
  assign new_n2461_ = ((~P1_EBX_REG_5__SCAN_IN | (new_n2091_ ? new_n2073_ : new_n2067_)) & (~P1_INSTADDRPOINTER_REG_5__SCAN_IN | (~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_))) ? (new_n2067_ | new_n2091_ | (P1_INSTADDRPOINTER_REG_4__SCAN_IN & (new_n2067_ | new_n2073_) & (new_n2073_ | ~new_n2116_)) | (P1_EBX_REG_4__SCAN_IN & (new_n2091_ ? ~new_n2073_ : ~new_n2067_))) : ((~new_n2067_ & ~new_n2091_) | ((~P1_INSTADDRPOINTER_REG_4__SCAN_IN | (~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_)) & (~P1_EBX_REG_4__SCAN_IN | (new_n2091_ ? new_n2073_ : new_n2067_))));
  assign new_n2462_ = ((~P1_EBX_REG_7__SCAN_IN | (new_n2091_ ? new_n2073_ : new_n2067_)) & (~P1_INSTADDRPOINTER_REG_7__SCAN_IN | (~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_))) ? (new_n2067_ | new_n2091_ | (P1_INSTADDRPOINTER_REG_6__SCAN_IN & (new_n2067_ | new_n2073_) & (new_n2073_ | ~new_n2116_)) | (P1_EBX_REG_6__SCAN_IN & (new_n2091_ ? ~new_n2073_ : ~new_n2067_))) : ((~new_n2067_ & ~new_n2091_) | ((~P1_INSTADDRPOINTER_REG_6__SCAN_IN | (~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_)) & (~P1_EBX_REG_6__SCAN_IN | (new_n2091_ ? new_n2073_ : new_n2067_))));
  assign new_n2463_ = ~new_n2465_ & (~new_n2464_ | (new_n2090_ & (new_n2455_ | ~P1_EBX_REG_8__SCAN_IN) & (~new_n2456_ | ~P1_INSTADDRPOINTER_REG_8__SCAN_IN))) & ~new_n2466_ & (new_n2464_ | (~new_n2090_ & ((~new_n2455_ & P1_EBX_REG_8__SCAN_IN) | (new_n2456_ & P1_INSTADDRPOINTER_REG_8__SCAN_IN))));
  assign new_n2464_ = (~P1_EBX_REG_9__SCAN_IN | (new_n2091_ ? new_n2073_ : new_n2067_)) & (~P1_INSTADDRPOINTER_REG_9__SCAN_IN | (~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_));
  assign new_n2465_ = (~P1_EBX_REG_11__SCAN_IN | (new_n2091_ ? new_n2073_ : new_n2067_)) & (~P1_INSTADDRPOINTER_REG_11__SCAN_IN | (~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_)) & ((P1_INSTADDRPOINTER_REG_10__SCAN_IN & (new_n2067_ | new_n2073_) & (new_n2073_ | ~new_n2116_)) | (P1_EBX_REG_10__SCAN_IN & (new_n2091_ ? ~new_n2073_ : ~new_n2067_)));
  assign new_n2466_ = (~new_n2067_ & ~new_n2091_) ? ((P1_EBX_REG_11__SCAN_IN & (new_n2091_ ? ~new_n2073_ : ~new_n2067_)) | (P1_INSTADDRPOINTER_REG_11__SCAN_IN & (new_n2067_ | new_n2073_) & (new_n2073_ | ~new_n2116_))) : ((~P1_INSTADDRPOINTER_REG_10__SCAN_IN | (~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_)) & (~P1_EBX_REG_10__SCAN_IN | (new_n2091_ ? new_n2073_ : new_n2067_)));
  assign new_n2467_ = ~new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_12__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_12__SCAN_IN));
  assign new_n2468_ = ~new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_13__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_13__SCAN_IN));
  assign new_n2469_ = ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_15__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_15__SCAN_IN)) ? (~new_n2090_ | (~new_n2455_ & P1_EBX_REG_14__SCAN_IN) | (new_n2456_ & P1_INSTADDRPOINTER_REG_14__SCAN_IN)) : (new_n2090_ | ((new_n2455_ | ~P1_EBX_REG_14__SCAN_IN) & (~new_n2456_ | ~P1_INSTADDRPOINTER_REG_14__SCAN_IN)));
  assign new_n2470_ = ~new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_17__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_17__SCAN_IN));
  assign new_n2471_ = ~new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_18__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_18__SCAN_IN));
  assign new_n2472_ = ~new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_22__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_22__SCAN_IN));
  assign new_n2473_ = ~new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_19__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_19__SCAN_IN));
  assign new_n2474_ = ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_21__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_21__SCAN_IN)) ? (~new_n2090_ | (~new_n2455_ & P1_EBX_REG_20__SCAN_IN) | (new_n2456_ & P1_INSTADDRPOINTER_REG_20__SCAN_IN)) : (new_n2090_ | ((new_n2455_ | ~P1_EBX_REG_20__SCAN_IN) & (~new_n2456_ | ~P1_INSTADDRPOINTER_REG_20__SCAN_IN)));
  assign new_n2475_ = ~new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_23__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_23__SCAN_IN));
  assign new_n2476_ = new_n2495_ & ((new_n2106_ & new_n2494_) | (new_n2477_ & new_n2493_));
  assign new_n2477_ = ~new_n2478_ & ~new_n2482_;
  assign new_n2478_ = new_n2479_ & new_n2136_ & (~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN) & (new_n2480_ | (~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN));
  assign new_n2479_ = ~new_n2065_ & ~new_n2067_;
  assign new_n2480_ = (~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & ((~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) | ((~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & ((~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN) | ((~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (new_n2481_ | (~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN))))));
  assign new_n2481_ = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign new_n2482_ = ~new_n2492_ & (~new_n2491_ | (new_n2489_ & ((~new_n2483_ & ~new_n2486_ & (~new_n2484_ | new_n2485_)) | new_n2487_ | (~new_n2484_ & new_n2485_))));
  assign new_n2483_ = ~new_n2065_ & ~new_n2067_ & ~new_n2079_ & ~new_n2073_ & P1_STATE2_REG_0__SCAN_IN & ((~new_n2073_ & P1_STATE2_REG_0__SCAN_IN & (new_n2079_ ? ~new_n2065_ : (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ^ ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN))) | (P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN) | ((~new_n2065_ | new_n2073_) & new_n2067_ & P1_STATE2_REG_0__SCAN_IN) | ((~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & P1_STATE2_REG_0__SCAN_IN & (new_n2073_ | new_n2079_)));
  assign new_n2484_ = P1_STATE2_REG_0__SCAN_IN & ((~new_n2073_ & ~new_n2079_ & ~new_n2065_ & ~new_n2067_) | (new_n2481_ ^ (P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN)));
  assign new_n2485_ = ((new_n2481_ ^ (P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN)) | new_n2079_ | new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN) & (~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_STATE2_REG_0__SCAN_IN) & (~new_n2065_ | ~P1_STATE2_REG_0__SCAN_IN) & (new_n2067_ | ~new_n2079_ | ~P1_STATE2_REG_0__SCAN_IN) & (~P1_STATE2_REG_0__SCAN_IN | new_n2067_ | ~new_n2073_);
  assign new_n2486_ = ((~new_n2073_ & P1_STATE2_REG_0__SCAN_IN & (new_n2079_ ? ~new_n2065_ : (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ^ ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN))) | (P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN) | ((~new_n2065_ | new_n2073_) & new_n2067_ & P1_STATE2_REG_0__SCAN_IN)) & (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & P1_STATE2_REG_0__SCAN_IN & (new_n2073_ | new_n2079_);
  assign new_n2487_ = (~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_STATE2_REG_0__SCAN_IN) & ((new_n2065_ & ~new_n2073_) | ~new_n2067_ | ~P1_STATE2_REG_0__SCAN_IN) & (~new_n2488_ | ~P1_STATE2_REG_0__SCAN_IN | (~new_n2073_ & ~new_n2079_)) & (new_n2488_ | new_n2079_ | new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN);
  assign new_n2488_ = ((~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (new_n2481_ | (~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN))) ^ (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2489_ = (~new_n2488_ | ~P1_STATE2_REG_0__SCAN_IN | (~new_n2073_ & ~new_n2079_) | ((~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_STATE2_REG_0__SCAN_IN) & ((new_n2065_ & ~new_n2073_) | ~new_n2067_ | ~P1_STATE2_REG_0__SCAN_IN))) & (new_n2073_ | new_n2079_ | new_n2065_ | new_n2067_ | new_n2490_ | ~P1_STATE2_REG_0__SCAN_IN);
  assign new_n2490_ = ((~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & ((~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN) | ((~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (new_n2481_ | (~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN))))) ^ (P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ^ ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n2491_ = (P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_STATE2_REG_0__SCAN_IN) & (~P1_STATE2_REG_0__SCAN_IN | (~new_n2073_ & ~new_n2079_) | (new_n2490_ & (~new_n2480_ | (~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN)) & (new_n2480_ | (~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ^ P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN))));
  assign new_n2492_ = (P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P1_STATE2_REG_0__SCAN_IN) & ((~new_n2073_ & ~new_n2079_ & ~new_n2065_ & ~new_n2067_ & (~new_n2480_ ^ (P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ^ ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN))) | ~P1_STATE2_REG_0__SCAN_IN | ((new_n2073_ | new_n2079_) & (~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN) & (new_n2480_ | (~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN))));
  assign new_n2493_ = ~new_n2073_ & ~new_n2091_ & ~new_n2067_ & new_n2097_ & ~new_n2065_ & ~new_n2053_ & ~new_n2079_ & new_n2085_;
  assign new_n2494_ = ~new_n2067_ & ~new_n2073_;
  assign new_n2495_ = new_n2118_ & P1_STATE2_REG_0__SCAN_IN;
  assign new_n2496_ = (((new_n2455_ | ~P1_EBX_REG_27__SCAN_IN) & (~new_n2456_ | ~P1_INSTADDRPOINTER_REG_27__SCAN_IN)) | (~new_n2090_ & ((new_n2456_ & P1_INSTADDRPOINTER_REG_26__SCAN_IN) | (~new_n2455_ & P1_EBX_REG_26__SCAN_IN)))) & (new_n2497_ | (~new_n2455_ & P1_EBX_REG_27__SCAN_IN) | (new_n2456_ & P1_INSTADDRPOINTER_REG_27__SCAN_IN)) & (~new_n2497_ | (new_n2090_ & (~new_n2456_ | ~P1_INSTADDRPOINTER_REG_26__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_26__SCAN_IN)));
  assign new_n2497_ = (~new_n2456_ | ~P1_INSTADDRPOINTER_REG_28__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_28__SCAN_IN);
  assign new_n2498_ = ~new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_29__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_29__SCAN_IN));
  assign new_n2499_ = ~new_n2500_ & ~new_n2514_ & new_n2518_ & ~new_n2608_ & new_n4452_ & ~new_n4467_ & new_n2623_ & new_n2654_;
  assign new_n2500_ = (new_n2503_ | new_n2504_) & (~new_n2501_ | new_n2502_) & (new_n2501_ | ~new_n2502_);
  assign new_n2501_ = (~new_n2324_ | ~new_n2425_) & ((~new_n2324_ & ~new_n2425_) | ((~new_n2324_ | ~new_n2432_) & ((~new_n2324_ & ~new_n2432_) | (~new_n2044_ & new_n2422_))));
  assign new_n2502_ = new_n2324_ ^ new_n2369_;
  assign new_n2503_ = new_n2476_ & ~new_n2053_;
  assign new_n2504_ = new_n2505_ & new_n2512_;
  assign new_n2505_ = new_n2118_ & (new_n2506_ | (new_n2106_ & new_n2111_) | (new_n2511_ & ~new_n2477_ & P1_STATE2_REG_0__SCAN_IN));
  assign new_n2506_ = ~new_n2510_ & (new_n2507_ | ((new_n2478_ | new_n2482_) & P1_STATE2_REG_0__SCAN_IN & new_n2494_ & new_n2509_));
  assign new_n2507_ = new_n2129_ & new_n2508_;
  assign new_n2508_ = ((P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (~new_n2480_ & (P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN))) & (~new_n2490_ | (new_n2480_ & (P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN) & (~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN)) | (~new_n2480_ & (P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ^ P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN)) | ~new_n2488_ | (new_n2481_ & (P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN)) | (~new_n2481_ & (P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN)));
  assign new_n2509_ = new_n2065_ & new_n2079_ & ~new_n2053_ & new_n2085_ & new_n2097_ & ~new_n2091_;
  assign new_n2510_ = READY1 & READY11_REG_SCAN_IN;
  assign new_n2511_ = ~new_n2091_ & new_n2067_ & new_n2073_ & new_n2097_ & ~new_n2065_ & ~new_n2053_ & ~new_n2079_ & new_n2085_;
  assign new_n2512_ = ~new_n2291_ & ~new_n2513_;
  assign new_n2513_ = ~new_n2053_ & new_n2065_;
  assign new_n2514_ = (~new_n2476_ | new_n2053_ | (new_n2515_ & ~new_n2516_) | (~new_n2515_ & new_n2516_)) & (new_n2476_ | ~P1_EBX_REG_22__SCAN_IN) & (~new_n2517_ | ~new_n2476_ | ~new_n2053_);
  assign new_n2515_ = (~new_n2324_ | ~new_n2432_) & ((~new_n2324_ & ~new_n2432_) | (~new_n2044_ & new_n2422_));
  assign new_n2516_ = new_n2324_ ^ new_n2425_;
  assign new_n2517_ = new_n2472_ ^ (~new_n2474_ & new_n2453_ & new_n2473_);
  assign new_n2518_ = new_n2600_ & ~new_n2520_ & ((~new_n2519_ & (new_n1929_ | P2_INSTADDRPOINTER_REG_17__SCAN_IN) & (~new_n1929_ | ~P2_INSTADDRPOINTER_REG_17__SCAN_IN)) | ~new_n2040_ | (new_n2519_ & (new_n1929_ ^ ~P2_INSTADDRPOINTER_REG_17__SCAN_IN)));
  assign new_n2519_ = (~new_n1922_ | ~P2_INSTADDRPOINTER_REG_16__SCAN_IN) & ((~new_n1922_ & ~P2_INSTADDRPOINTER_REG_16__SCAN_IN) | (new_n1936_ & (~new_n1933_ | new_n1930_ | (~new_n1932_ & (new_n1797_ | new_n1927_)))));
  assign new_n2520_ = new_n2562_ & ((P1_INSTADDRPOINTER_REG_24__SCAN_IN & ((~new_n2561_ & (~new_n2521_ | ~new_n2560_)) | (~new_n2558_ & P1_INSTADDRPOINTER_REG_23__SCAN_IN)) & ((new_n2521_ & new_n2560_) | (new_n2558_ & ~P1_INSTADDRPOINTER_REG_23__SCAN_IN))) | ~new_n2596_ | (~P1_INSTADDRPOINTER_REG_24__SCAN_IN & (((new_n2561_ | (new_n2521_ & new_n2560_)) & (new_n2558_ | ~P1_INSTADDRPOINTER_REG_23__SCAN_IN)) | ((~new_n2521_ | ~new_n2560_) & (~new_n2558_ | P1_INSTADDRPOINTER_REG_23__SCAN_IN)))));
  assign new_n2521_ = new_n2559_ & (~new_n2557_ | (~new_n2555_ & (new_n2522_ | ~new_n2552_)));
  assign new_n2522_ = ~new_n2550_ & new_n2551_ & ~new_n2549_ & (new_n2523_ | (new_n2548_ & (~new_n2546_ | (~new_n2524_ & ~new_n2530_))));
  assign new_n2523_ = P1_INSTADDRPOINTER_REG_11__SCAN_IN & new_n2479_ & (~new_n2305_ | new_n2202_) & (new_n2305_ | ~new_n2202_);
  assign new_n2524_ = new_n2525_ & ~P1_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign new_n2525_ = (~new_n2479_ | (new_n2048_ & new_n2221_) | (~new_n2048_ & ~new_n2221_)) & (~new_n2529_ | new_n2164_ | ~new_n2526_ | new_n2179_);
  assign new_n2526_ = new_n2527_ & ~new_n2186_;
  assign new_n2527_ = ~new_n2193_ & ~new_n2138_ & (new_n2528_ | ~new_n2149_);
  assign new_n2528_ = ~new_n2170_ & ~new_n2158_;
  assign new_n2529_ = new_n2067_ & ~new_n2073_;
  assign new_n2530_ = (new_n2531_ | ~P1_INSTADDRPOINTER_REG_7__SCAN_IN) & ((new_n2531_ & ~P1_INSTADDRPOINTER_REG_7__SCAN_IN) | ((new_n2533_ | ~P1_INSTADDRPOINTER_REG_6__SCAN_IN) & ((new_n2533_ & ~P1_INSTADDRPOINTER_REG_6__SCAN_IN) | ((new_n2534_ | ~P1_INSTADDRPOINTER_REG_5__SCAN_IN) & (new_n2535_ | (new_n2534_ & ~P1_INSTADDRPOINTER_REG_5__SCAN_IN))))));
  assign new_n2531_ = ~new_n2532_ & (~new_n2479_ | (new_n2252_ & (~new_n2251_ | new_n2198_)) | new_n2255_ | (new_n2253_ & (new_n2251_ | new_n2185_)));
  assign new_n2532_ = (~new_n2164_ | (new_n2526_ & ~new_n2179_)) & new_n2529_ & (new_n2164_ | ~new_n2526_ | new_n2179_);
  assign new_n2533_ = (~new_n2479_ | (new_n2257_ & (new_n2198_ | (~new_n2251_ & ~new_n2185_))) | (~new_n2257_ & ~new_n2198_ & (new_n2251_ | new_n2185_))) & ((~new_n2526_ & new_n2179_) | ~new_n2529_ | (new_n2526_ & ~new_n2179_));
  assign new_n2534_ = (~new_n2261_ | ~new_n2479_) & ((~new_n2527_ & new_n2186_) | ~new_n2529_ | (new_n2527_ & ~new_n2186_));
  assign new_n2535_ = (new_n2536_ | ~P1_INSTADDRPOINTER_REG_4__SCAN_IN) & ((new_n2536_ & ~P1_INSTADDRPOINTER_REG_4__SCAN_IN) | ((new_n2538_ | ~P1_INSTADDRPOINTER_REG_3__SCAN_IN) & ((new_n2538_ & ~P1_INSTADDRPOINTER_REG_3__SCAN_IN) | ((new_n2540_ | ~P1_INSTADDRPOINTER_REG_2__SCAN_IN) & (~new_n2542_ | (new_n2540_ & ~P1_INSTADDRPOINTER_REG_2__SCAN_IN))))));
  assign new_n2536_ = ~new_n2537_ & (~new_n2479_ | (new_n2270_ ^ (~new_n2049_ & (new_n2147_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))))));
  assign new_n2537_ = (~new_n2193_ | (~new_n2138_ & (new_n2528_ | ~new_n2149_))) & new_n2529_ & (new_n2193_ | new_n2138_ | (~new_n2528_ & new_n2149_));
  assign new_n2538_ = (~new_n2479_ | (~new_n2277_ & (new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_))) | (new_n2277_ & ((~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))))) & ((new_n2539_ & new_n2138_) | ~new_n2529_ | (~new_n2539_ & ~new_n2138_));
  assign new_n2539_ = ~new_n2528_ & new_n2149_;
  assign new_n2540_ = (~new_n2479_ | (new_n2154_ & ~new_n2283_) | (~new_n2154_ & new_n2283_)) & ~new_n2541_ & (~new_n2529_ | (new_n2528_ ^ ~new_n2149_));
  assign new_n2541_ = new_n2073_ & ~new_n2091_;
  assign new_n2542_ = (P1_INSTADDRPOINTER_REG_1__SCAN_IN | (~new_n2543_ & P1_INSTADDRPOINTER_REG_0__SCAN_IN)) & ((new_n2284_ & new_n2479_) | ~new_n2544_ | (~new_n2543_ & P1_INSTADDRPOINTER_REG_1__SCAN_IN & P1_INSTADDRPOINTER_REG_0__SCAN_IN));
  assign new_n2543_ = (~new_n2479_ | (new_n2156_ & ~new_n2288_) | (~new_n2156_ & new_n2288_)) & ~new_n2541_ & (~new_n2529_ | ~new_n2158_);
  assign new_n2544_ = ((new_n2170_ & new_n2158_) | ~new_n2067_ | new_n2073_ | (~new_n2170_ & ~new_n2158_)) & new_n2545_ & (~new_n2065_ | new_n2073_);
  assign new_n2545_ = new_n2097_ & ~new_n2091_;
  assign new_n2546_ = (~P1_INSTADDRPOINTER_REG_10__SCAN_IN | ~new_n2306_ | ~new_n2479_) & (new_n2525_ | ~P1_INSTADDRPOINTER_REG_8__SCAN_IN) & (~new_n2547_ | ~P1_INSTADDRPOINTER_REG_9__SCAN_IN);
  assign new_n2547_ = new_n2479_ & (new_n2215_ | new_n2048_ | new_n2221_) & (~new_n2215_ | (~new_n2048_ & ~new_n2221_));
  assign new_n2548_ = (new_n2547_ | P1_INSTADDRPOINTER_REG_9__SCAN_IN | (P1_INSTADDRPOINTER_REG_10__SCAN_IN & new_n2306_ & new_n2479_)) & (P1_INSTADDRPOINTER_REG_10__SCAN_IN | (new_n2306_ & new_n2479_)) & (P1_INSTADDRPOINTER_REG_11__SCAN_IN | (new_n2479_ & (new_n2305_ | ~new_n2202_) & (~new_n2305_ | new_n2202_)));
  assign new_n2549_ = ~P1_INSTADDRPOINTER_REG_12__SCAN_IN & (~new_n2479_ | (new_n2047_ & ~new_n2244_) | (~new_n2047_ & new_n2244_));
  assign new_n2550_ = ~P1_INSTADDRPOINTER_REG_13__SCAN_IN & (~new_n2479_ | ((~new_n2227_ ^ ~new_n2163_) & new_n2047_ & (new_n2232_ ^ new_n2163_)) | ((~new_n2227_ | new_n2163_) & (new_n2227_ | ~new_n2163_) & (~new_n2047_ | (~new_n2232_ ^ new_n2163_))));
  assign new_n2551_ = (P1_INSTADDRPOINTER_REG_14__SCAN_IN | (new_n2479_ & (~new_n2309_ | (new_n2311_ ^ ~new_n2163_)) & (new_n2309_ | (new_n2311_ & ~new_n2163_) | (~new_n2311_ & new_n2163_)))) & (P1_INSTADDRPOINTER_REG_15__SCAN_IN | (new_n2479_ & ((~new_n2316_ ^ new_n2163_) | ~new_n2309_ | (new_n2311_ ^ ~new_n2163_)) & ((~new_n2316_ & new_n2163_) | (new_n2316_ & ~new_n2163_) | (new_n2309_ & (~new_n2311_ ^ ~new_n2163_)))));
  assign new_n2552_ = (~P1_INSTADDRPOINTER_REG_15__SCAN_IN | ~new_n2479_ | (~new_n2554_ & new_n2309_ & ~new_n2326_) | (new_n2554_ & (~new_n2309_ | new_n2326_))) & ((~P1_INSTADDRPOINTER_REG_14__SCAN_IN & (~new_n2479_ | (~new_n2309_ & new_n2326_) | (new_n2309_ & ~new_n2326_))) | (~P1_INSTADDRPOINTER_REG_15__SCAN_IN & (~new_n2479_ | (~new_n2554_ & new_n2309_ & ~new_n2326_) | (new_n2554_ & (~new_n2309_ | new_n2326_)))) | (new_n2553_ & (~P1_INSTADDRPOINTER_REG_14__SCAN_IN | ~new_n2479_ | (~new_n2309_ & new_n2326_) | (new_n2309_ & ~new_n2326_))));
  assign new_n2553_ = (~P1_INSTADDRPOINTER_REG_13__SCAN_IN | ~new_n2479_ | ((~new_n2227_ ^ ~new_n2163_) & new_n2047_ & (new_n2232_ ^ new_n2163_)) | ((~new_n2227_ | new_n2163_) & (new_n2227_ | ~new_n2163_) & (~new_n2047_ | (~new_n2232_ ^ new_n2163_)))) & ((~P1_INSTADDRPOINTER_REG_13__SCAN_IN & (~new_n2479_ | ((~new_n2227_ ^ ~new_n2163_) & new_n2047_ & (new_n2232_ ^ new_n2163_)) | ((~new_n2227_ | new_n2163_) & (new_n2227_ | ~new_n2163_) & (~new_n2047_ | (~new_n2232_ ^ new_n2163_))))) | ~P1_INSTADDRPOINTER_REG_12__SCAN_IN | ~new_n2479_ | (new_n2047_ & (new_n2232_ ^ new_n2163_)) | (~new_n2047_ & (new_n2232_ | ~new_n2163_) & (~new_n2232_ | new_n2163_)));
  assign new_n2554_ = new_n2316_ ^ ~new_n2163_;
  assign new_n2555_ = ~new_n2556_ & ~P1_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign new_n2556_ = new_n2479_ & ((new_n2163_ & (~new_n2325_ | (~new_n2316_ ^ new_n2163_))) | (new_n2325_ & new_n2316_ & ~new_n2163_));
  assign new_n2557_ = (~new_n2556_ | ~P1_INSTADDRPOINTER_REG_16__SCAN_IN) & (~new_n2558_ | ~P1_INSTADDRPOINTER_REG_17__SCAN_IN);
  assign new_n2558_ = new_n2479_ & new_n2163_ & (~new_n2325_ | (~new_n2316_ ^ new_n2163_));
  assign new_n2559_ = (new_n2558_ | P1_INSTADDRPOINTER_REG_17__SCAN_IN) & (new_n2558_ | P1_INSTADDRPOINTER_REG_18__SCAN_IN);
  assign new_n2560_ = (new_n2558_ | (P1_INSTADDRPOINTER_REG_22__SCAN_IN & P1_INSTADDRPOINTER_REG_21__SCAN_IN)) & (new_n2558_ | P1_INSTADDRPOINTER_REG_20__SCAN_IN) & (new_n2558_ | P1_INSTADDRPOINTER_REG_19__SCAN_IN);
  assign new_n2561_ = new_n2558_ & (P1_INSTADDRPOINTER_REG_22__SCAN_IN | P1_INSTADDRPOINTER_REG_18__SCAN_IN | P1_INSTADDRPOINTER_REG_21__SCAN_IN | P1_INSTADDRPOINTER_REG_20__SCAN_IN | P1_INSTADDRPOINTER_REG_19__SCAN_IN);
  assign new_n2562_ = ~new_n2563_ & ~new_n2573_ & (~new_n2588_ | (new_n2590_ & P1_INSTADDRPOINTER_REG_24__SCAN_IN) | (~new_n2590_ & ~P1_INSTADDRPOINTER_REG_24__SCAN_IN)) & (~new_n2589_ | ~P1_REIP_REG_24__SCAN_IN);
  assign new_n2563_ = (new_n2452_ | (~new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_24__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_24__SCAN_IN)))) & new_n2564_ & (~new_n2452_ | (~new_n2090_ & (~new_n2456_ | ~P1_INSTADDRPOINTER_REG_24__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_24__SCAN_IN)) | (new_n2090_ & ((new_n2456_ & P1_INSTADDRPOINTER_REG_24__SCAN_IN) | (~new_n2455_ & P1_EBX_REG_24__SCAN_IN))));
  assign new_n2564_ = new_n2565_ & ~new_n2572_;
  assign new_n2565_ = new_n2495_ & (new_n2566_ | ~new_n2568_);
  assign new_n2566_ = (new_n2067_ | (new_n2567_ & (new_n2478_ | new_n2482_))) & ~new_n2097_ & ~new_n2510_ & (new_n2508_ | ~new_n2067_);
  assign new_n2567_ = ~new_n2116_ & ~P1_STATE_REG_0__SCAN_IN;
  assign new_n2568_ = (~new_n2569_ | (~new_n2478_ & ~new_n2482_)) & new_n2571_ & (new_n2478_ | new_n2482_ | ~new_n2570_ | new_n2067_);
  assign new_n2569_ = new_n2097_ & (new_n2291_ | new_n2073_ | (new_n2509_ & ~new_n2510_ & (~new_n2067_ | new_n2567_)));
  assign new_n2570_ = new_n2097_ & ~new_n2065_ & ~new_n2053_ & ~new_n2079_ & new_n2085_;
  assign new_n2571_ = (~new_n2097_ | ((~new_n2073_ | (~new_n2065_ & ~new_n2053_ & ~new_n2079_ & new_n2085_)) & ~new_n2091_ & ~new_n2053_ & (~new_n2065_ | new_n2085_) & (~new_n2085_ | new_n2065_ | ~new_n2079_))) & (new_n2097_ | (new_n2073_ & new_n2091_ & ~new_n2065_ & new_n2079_ & ~new_n2053_ & ~new_n2085_)) & (~new_n2067_ | new_n2073_ | ((~new_n2065_ | new_n2085_) & ((~new_n2053_ & new_n2065_) | (~new_n2053_ & ~new_n2085_)))) & (new_n2073_ | new_n2079_ | (~new_n2065_ & new_n2085_));
  assign new_n2572_ = (~new_n2529_ | ~new_n2509_) & (~new_n2096_ | ~new_n2079_);
  assign new_n2573_ = (P1_INSTADDRPOINTER_REG_24__SCAN_IN | (new_n2577_ & P1_INSTADDRPOINTER_REG_23__SCAN_IN & (new_n2584_ | (new_n2586_ & P1_INSTADDRPOINTER_REG_0__SCAN_IN)))) & (new_n2574_ | (new_n2586_ & (~P1_INSTADDRPOINTER_REG_23__SCAN_IN | ~new_n2577_ | ~P1_INSTADDRPOINTER_REG_0__SCAN_IN)) | ~P1_INSTADDRPOINTER_REG_24__SCAN_IN | (new_n2584_ & (~new_n2577_ | ~P1_INSTADDRPOINTER_REG_23__SCAN_IN)));
  assign new_n2574_ = ~new_n2565_ & ~new_n2575_;
  assign new_n2575_ = ~P1_STATE2_REG_0__SCAN_IN & new_n2576_ & ~P1_STATE2_REG_1__SCAN_IN;
  assign new_n2576_ = ~P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_2__SCAN_IN;
  assign new_n2577_ = P1_INSTADDRPOINTER_REG_22__SCAN_IN & P1_INSTADDRPOINTER_REG_21__SCAN_IN & P1_INSTADDRPOINTER_REG_20__SCAN_IN & new_n2583_ & new_n2578_ & P1_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign new_n2578_ = P1_INSTADDRPOINTER_REG_16__SCAN_IN & P1_INSTADDRPOINTER_REG_15__SCAN_IN & new_n2579_ & P1_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign new_n2579_ = new_n2580_ & P1_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign new_n2580_ = new_n2581_ & P1_INSTADDRPOINTER_REG_12__SCAN_IN & P1_INSTADDRPOINTER_REG_11__SCAN_IN & P1_INSTADDRPOINTER_REG_8__SCAN_IN & P1_INSTADDRPOINTER_REG_10__SCAN_IN & P1_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign new_n2581_ = P1_INSTADDRPOINTER_REG_7__SCAN_IN & new_n2582_ & P1_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign new_n2582_ = P1_INSTADDRPOINTER_REG_2__SCAN_IN & P1_INSTADDRPOINTER_REG_1__SCAN_IN & P1_INSTADDRPOINTER_REG_3__SCAN_IN & P1_INSTADDRPOINTER_REG_5__SCAN_IN & P1_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign new_n2583_ = P1_INSTADDRPOINTER_REG_19__SCAN_IN & P1_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign new_n2584_ = new_n2585_ & new_n2495_ & (new_n2566_ | ~new_n2568_);
  assign new_n2585_ = ~new_n2067_ & new_n2073_ & ~new_n2097_ & new_n2091_ & ~new_n2065_ & new_n2079_ & ~new_n2053_ & ~new_n2085_;
  assign new_n2586_ = ~new_n2587_ & new_n2495_ & (new_n2566_ | ~new_n2568_);
  assign new_n2587_ = ((new_n2067_ & (new_n2091_ | (~new_n2065_ & ~new_n2053_ & ~new_n2079_ & new_n2085_)) & (~new_n2053_ | (new_n2065_ & new_n2079_)) & ((new_n2065_ & ~new_n2085_) | ~new_n2097_ | (~new_n2079_ & new_n2085_)) & (new_n2097_ | ((~new_n2065_ | new_n2085_) & new_n2079_ & (new_n2053_ | ~new_n2085_)))) | ~new_n2073_ | (new_n2079_ & ~new_n2065_ & ~new_n2067_)) & (new_n2067_ | ((new_n2091_ | (~new_n2053_ & (~new_n2065_ | new_n2085_) & (~new_n2085_ | new_n2065_ | ~new_n2079_))) & (new_n2097_ | ~new_n2085_) & (~new_n2073_ | ~new_n2097_ | ~new_n2091_))) & (~new_n2067_ | new_n2073_ | ((~new_n2065_ | new_n2085_) & ((~new_n2053_ & new_n2065_) | (~new_n2053_ & ~new_n2085_)))) & (new_n2073_ | new_n2079_ | (~new_n2065_ & new_n2085_)) & ((new_n2097_ & ~new_n2091_) | (new_n2073_ & (new_n2067_ | new_n2091_))) & (~new_n2053_ | new_n2067_) & (~new_n2073_ | ~new_n2097_ | ~new_n2091_ | new_n2085_ | ~new_n2065_ | ~new_n2053_ | ~new_n2079_) & (~new_n2073_ | new_n2067_ | new_n2091_ | new_n2065_ | ~new_n2079_ | new_n2053_ | new_n2085_) & (new_n2097_ | ~new_n2085_ | ~new_n2065_ | ~new_n2053_ | ~new_n2079_) & (~new_n2067_ | ~new_n2073_ | ~new_n2097_ | ~new_n2091_ | new_n2053_ | new_n2079_ | ~new_n2085_);
  assign new_n2588_ = new_n2565_ & new_n2493_;
  assign new_n2589_ = ~P1_STATE2_REG_2__SCAN_IN & (new_n2575_ | (new_n2495_ & (new_n2566_ | ~new_n2568_)));
  assign new_n2590_ = new_n2591_ & P1_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign new_n2591_ = P1_INSTADDRPOINTER_REG_22__SCAN_IN & P1_INSTADDRPOINTER_REG_21__SCAN_IN & P1_INSTADDRPOINTER_REG_20__SCAN_IN & new_n2583_ & new_n2592_ & P1_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign new_n2592_ = P1_INSTADDRPOINTER_REG_16__SCAN_IN & P1_INSTADDRPOINTER_REG_15__SCAN_IN & new_n2593_ & P1_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign new_n2593_ = P1_INSTADDRPOINTER_REG_13__SCAN_IN & new_n2594_ & P1_INSTADDRPOINTER_REG_12__SCAN_IN & P1_INSTADDRPOINTER_REG_11__SCAN_IN & P1_INSTADDRPOINTER_REG_8__SCAN_IN & P1_INSTADDRPOINTER_REG_10__SCAN_IN & P1_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign new_n2594_ = P1_INSTADDRPOINTER_REG_7__SCAN_IN & new_n2595_ & P1_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign new_n2595_ = P1_INSTADDRPOINTER_REG_3__SCAN_IN & P1_INSTADDRPOINTER_REG_5__SCAN_IN & P1_INSTADDRPOINTER_REG_4__SCAN_IN & (P1_INSTADDRPOINTER_REG_2__SCAN_IN | (P1_INSTADDRPOINTER_REG_1__SCAN_IN & P1_INSTADDRPOINTER_REG_0__SCAN_IN));
  assign new_n2596_ = new_n2565_ & (new_n2511_ | ~new_n2597_ | new_n2599_ | (new_n2096_ & ~new_n2079_));
  assign new_n2597_ = (~P1_STATE2_REG_2__SCAN_IN | ~new_n2509_ | new_n2067_ | new_n2073_) & (~new_n2598_ | ~new_n2545_ | new_n2073_);
  assign new_n2598_ = ~new_n2065_ & new_n2079_ & ~new_n2053_ & ~new_n2085_;
  assign new_n2599_ = new_n2266_ & new_n2067_ & new_n2073_;
  assign new_n2600_ = (((new_n2044_ | (new_n2324_ & ~new_n2353_) | (new_n2324_ & new_n2360_)) & (new_n2324_ | new_n2432_) & (~new_n2324_ | ~new_n2432_)) | ~new_n2602_ | (~new_n2044_ & (~new_n2324_ | new_n2353_) & (~new_n2324_ | ~new_n2360_) & (new_n2324_ ^ ~new_n2432_))) & (((~new_n2324_ ^ ~new_n2353_) & ~new_n2601_ & (~new_n2324_ | ~new_n2360_)) | ~new_n2503_ | ((~new_n2324_ | new_n2353_) & (new_n2324_ | ~new_n2353_) & (new_n2601_ | (new_n2324_ & new_n2360_))));
  assign new_n2601_ = (new_n2324_ | new_n2360_) & ((new_n2324_ & new_n2346_) | ((new_n2324_ | new_n2346_) & ((new_n2324_ & ~new_n2339_) | ((new_n2324_ | ~new_n2339_) & (new_n2327_ | (~new_n2045_ & ~new_n2338_))))));
  assign new_n2602_ = ~new_n2603_ & P1_STATEBS16_REG_SCAN_IN & P1_STATE2_REG_1__SCAN_IN;
  assign new_n2603_ = ~new_n2604_ & ~new_n2606_;
  assign new_n2604_ = new_n2605_ & ~new_n2073_ & (new_n2478_ | new_n2482_);
  assign new_n2605_ = new_n2598_ & new_n2545_ & new_n2495_;
  assign new_n2606_ = ~new_n2607_ & ~P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN;
  assign new_n2607_ = P1_STATE2_REG_2__SCAN_IN & P1_STATE2_REG_1__SCAN_IN;
  assign new_n2608_ = ~new_n2609_ & new_n2618_ & ((~new_n2622_ & (~new_n2498_ | ~new_n2450_ | ~new_n2496_)) | ~new_n2564_ | (new_n2622_ & new_n2498_ & new_n2450_ & new_n2496_));
  assign new_n2609_ = (new_n2610_ | new_n2611_ | (~new_n2613_ & (new_n2616_ | (~new_n2614_ & new_n2521_ & new_n2560_)))) & new_n2596_ & (~new_n2610_ | (~new_n2611_ & (new_n2613_ | (~new_n2616_ & (new_n2614_ | ~new_n2521_ | ~new_n2560_)))));
  assign new_n2610_ = new_n2558_ ^ P1_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign new_n2611_ = new_n2558_ & (~new_n2612_ | P1_INSTADDRPOINTER_REG_29__SCAN_IN);
  assign new_n2612_ = ~P1_INSTADDRPOINTER_REG_24__SCAN_IN & ~P1_INSTADDRPOINTER_REG_23__SCAN_IN & ~P1_INSTADDRPOINTER_REG_26__SCAN_IN & ~P1_INSTADDRPOINTER_REG_25__SCAN_IN & ~P1_INSTADDRPOINTER_REG_21__SCAN_IN & ~P1_INSTADDRPOINTER_REG_20__SCAN_IN & ~P1_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign new_n2613_ = ~new_n2558_ & ~P1_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign new_n2614_ = ~new_n2558_ & ~new_n2615_;
  assign new_n2615_ = P1_INSTADDRPOINTER_REG_24__SCAN_IN & P1_INSTADDRPOINTER_REG_28__SCAN_IN & P1_INSTADDRPOINTER_REG_25__SCAN_IN & P1_INSTADDRPOINTER_REG_23__SCAN_IN & P1_INSTADDRPOINTER_REG_27__SCAN_IN & P1_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign new_n2616_ = new_n2558_ & ~new_n2617_;
  assign new_n2617_ = ~P1_INSTADDRPOINTER_REG_22__SCAN_IN & ~P1_INSTADDRPOINTER_REG_18__SCAN_IN & ~P1_INSTADDRPOINTER_REG_28__SCAN_IN & ~P1_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign new_n2618_ = new_n2619_ & ((~new_n2584_ & ~new_n2586_) | ((~P1_INSTADDRPOINTER_REG_30__SCAN_IN | (new_n2621_ & (~new_n2586_ | P1_INSTADDRPOINTER_REG_0__SCAN_IN))) & ((~new_n2584_ & ~P1_INSTADDRPOINTER_REG_0__SCAN_IN) | ~new_n2621_ | P1_INSTADDRPOINTER_REG_30__SCAN_IN)));
  assign new_n2619_ = (~P1_REIP_REG_30__SCAN_IN | new_n2574_ | P1_STATE2_REG_2__SCAN_IN) & (~new_n2574_ | ~P1_INSTADDRPOINTER_REG_30__SCAN_IN) & (~new_n2588_ | (~new_n2620_ & ~P1_INSTADDRPOINTER_REG_30__SCAN_IN) | (new_n2620_ & P1_INSTADDRPOINTER_REG_30__SCAN_IN));
  assign new_n2620_ = new_n2590_ & P1_INSTADDRPOINTER_REG_24__SCAN_IN & P1_INSTADDRPOINTER_REG_28__SCAN_IN & P1_INSTADDRPOINTER_REG_25__SCAN_IN & P1_INSTADDRPOINTER_REG_29__SCAN_IN & P1_INSTADDRPOINTER_REG_27__SCAN_IN & P1_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign new_n2621_ = new_n2577_ & P1_INSTADDRPOINTER_REG_23__SCAN_IN & P1_INSTADDRPOINTER_REG_24__SCAN_IN & P1_INSTADDRPOINTER_REG_28__SCAN_IN & P1_INSTADDRPOINTER_REG_25__SCAN_IN & P1_INSTADDRPOINTER_REG_29__SCAN_IN & P1_INSTADDRPOINTER_REG_27__SCAN_IN & P1_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign new_n2622_ = ~new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_30__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_30__SCAN_IN));
  assign new_n2623_ = new_n2625_ & (new_n2624_ | ~new_n2650_ | ((P2_INSTADDRPOINTER_REG_14__SCAN_IN | (new_n1959_ & P2_INSTADDRPOINTER_REG_13__SCAN_IN)) & new_n2028_ & (~new_n1959_ | ~P2_INSTADDRPOINTER_REG_13__SCAN_IN | ~P2_INSTADDRPOINTER_REG_14__SCAN_IN)));
  assign new_n2624_ = ((new_n1935_ ^ P2_INSTADDRPOINTER_REG_14__SCAN_IN) | ((new_n1931_ | P2_INSTADDRPOINTER_REG_13__SCAN_IN) & ((~new_n1797_ & ~new_n1927_) | (new_n1931_ & P2_INSTADDRPOINTER_REG_13__SCAN_IN)))) & new_n2040_ & ((new_n1935_ & P2_INSTADDRPOINTER_REG_14__SCAN_IN) | (~new_n1935_ & ~P2_INSTADDRPOINTER_REG_14__SCAN_IN) | (~new_n1931_ & ~P2_INSTADDRPOINTER_REG_13__SCAN_IN) | ((new_n1797_ | new_n1927_) & (~new_n1931_ | ~P2_INSTADDRPOINTER_REG_13__SCAN_IN)));
  assign new_n2625_ = (~new_n2627_ | (new_n2649_ & (new_n2626_ | (new_n2324_ & new_n2346_) | (~new_n2324_ & ~new_n2346_)) & (~new_n2626_ | (new_n2324_ ^ new_n2346_)))) & (~new_n2648_ | (new_n2503_ & (new_n2626_ | (new_n2324_ & new_n2346_) | (~new_n2324_ & ~new_n2346_)) & (~new_n2626_ | (new_n2324_ ^ new_n2346_))));
  assign new_n2626_ = (~new_n2324_ | new_n2339_) & ((~new_n2324_ & new_n2339_) | (~new_n2327_ & (new_n2045_ | new_n2338_)));
  assign new_n2627_ = (~new_n2639_ | ~new_n2645_) & (~new_n2643_ | (new_n2347_ & P1_PHYADDRPOINTER_REG_18__SCAN_IN) | (~new_n2347_ & ~P1_PHYADDRPOINTER_REG_18__SCAN_IN)) & new_n2628_ & (new_n2640_ | ~P1_EBX_REG_18__SCAN_IN);
  assign new_n2628_ = new_n2635_ & (~new_n2629_ | (new_n2637_ & new_n2471_) | (~new_n2637_ & ~new_n2471_));
  assign new_n2629_ = P1_EBX_REG_31__SCAN_IN & ~new_n2634_ & ~new_n2630_ & new_n2494_ & P1_STATE2_REG_2__SCAN_IN;
  assign new_n2630_ = new_n2633_ & (~new_n2118_ | (~new_n2631_ & new_n2632_));
  assign new_n2631_ = new_n2509_ & new_n2495_ & ~new_n2073_ & (new_n2478_ | new_n2482_);
  assign new_n2632_ = ~new_n2507_ & (~new_n2585_ | ~P1_STATE2_REG_0__SCAN_IN | (~new_n2478_ & ~new_n2482_));
  assign new_n2633_ = (P1_STATE2_REG_0__SCAN_IN | P1_STATE2_REG_1__SCAN_IN | P1_STATE2_REG_3__SCAN_IN | P1_STATE2_REG_2__SCAN_IN) & (P1_STATEBS16_REG_SCAN_IN | P1_STATE2_REG_2__SCAN_IN | ~P1_STATE2_REG_1__SCAN_IN | P1_STATE2_REG_0__SCAN_IN) & (P1_STATE2_REG_2__SCAN_IN | P1_STATE2_REG_1__SCAN_IN | ~P1_STATE2_REG_3__SCAN_IN | ~P1_STATE2_REG_0__SCAN_IN);
  assign new_n2634_ = ~new_n2510_ & ~P1_STATEBS16_REG_SCAN_IN;
  assign new_n2635_ = ~new_n2636_ & (~new_n2630_ | ~P1_REIP_REG_18__SCAN_IN) & (~P1_PHYADDRPOINTER_REG_18__SCAN_IN | new_n2630_ | ~P1_STATE2_REG_3__SCAN_IN);
  assign new_n2636_ = ~P1_STATE2_REG_1__SCAN_IN & ~P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_2__SCAN_IN & (~new_n2633_ | (P1_STATE2_REG_2__SCAN_IN & ~P1_STATE2_REG_1__SCAN_IN & (new_n2631_ | ~new_n2632_)));
  assign new_n2637_ = new_n2470_ & new_n2454_ & ~new_n2469_ & new_n2638_ & new_n2468_;
  assign new_n2638_ = new_n2467_ & new_n2457_ & new_n2463_;
  assign new_n2639_ = new_n2634_ & ((~new_n2630_ & new_n2494_ & P1_STATE2_REG_2__SCAN_IN) | (new_n2567_ & new_n2529_ & ~new_n2630_ & P1_STATE2_REG_2__SCAN_IN));
  assign new_n2640_ = ~new_n2641_ & ~new_n2642_;
  assign new_n2641_ = ~P1_EBX_REG_31__SCAN_IN & ~new_n2634_ & new_n2494_ & P1_STATE2_REG_2__SCAN_IN & (~new_n2633_ | (P1_STATE2_REG_2__SCAN_IN & ~P1_STATE2_REG_1__SCAN_IN & (new_n2631_ | ~new_n2632_)));
  assign new_n2642_ = (~new_n2567_ | ~new_n2634_) & new_n2529_ & P1_STATE2_REG_2__SCAN_IN & (~new_n2633_ | (P1_STATE2_REG_2__SCAN_IN & ~P1_STATE2_REG_1__SCAN_IN & (new_n2631_ | ~new_n2632_)));
  assign new_n2643_ = new_n2644_ & new_n2275_ & P1_STATE2_REG_1__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN;
  assign new_n2644_ = ~P1_PHYADDRPOINTER_REG_31__SCAN_IN ^ (P1_PHYADDRPOINTER_REG_30__SCAN_IN & P1_PHYADDRPOINTER_REG_29__SCAN_IN & P1_PHYADDRPOINTER_REG_28__SCAN_IN & new_n2418_ & P1_PHYADDRPOINTER_REG_27__SCAN_IN);
  assign new_n2645_ = P1_REIP_REG_18__SCAN_IN ^ (P1_REIP_REG_15__SCAN_IN & P1_REIP_REG_17__SCAN_IN & P1_REIP_REG_16__SCAN_IN & P1_REIP_REG_14__SCAN_IN & new_n2646_ & P1_REIP_REG_13__SCAN_IN & P1_REIP_REG_12__SCAN_IN);
  assign new_n2646_ = new_n2647_ & P1_REIP_REG_6__SCAN_IN & P1_REIP_REG_11__SCAN_IN & P1_REIP_REG_10__SCAN_IN & P1_REIP_REG_7__SCAN_IN & P1_REIP_REG_9__SCAN_IN & P1_REIP_REG_8__SCAN_IN;
  assign new_n2647_ = P1_REIP_REG_3__SCAN_IN & P1_REIP_REG_2__SCAN_IN & P1_REIP_REG_1__SCAN_IN & P1_REIP_REG_5__SCAN_IN & P1_REIP_REG_4__SCAN_IN;
  assign new_n2648_ = (new_n2476_ | ~P1_EBX_REG_18__SCAN_IN) & (~new_n2476_ | ~new_n2053_ | (~new_n2637_ & ~new_n2471_) | (new_n2637_ & new_n2471_));
  assign new_n2649_ = ~new_n2644_ & new_n2275_ & P1_STATE2_REG_1__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN;
  assign new_n2650_ = new_n2652_ & ((~new_n2651_ & new_n1992_) | ~new_n2004_ | (new_n2651_ & ~new_n1992_));
  assign new_n2651_ = ~new_n1991_ & new_n1988_ & ~new_n1987_ & ~new_n1986_ & ~new_n1985_ & new_n1978_ & ~new_n1984_;
  assign new_n2652_ = (~new_n2005_ | ~P2_PHYADDRPOINTER_REG_14__SCAN_IN) & (~P2_REIP_REG_14__SCAN_IN | new_n2005_ | ~new_n2022_) & (new_n2005_ | new_n2021_ | (new_n2653_ & P2_PHYADDRPOINTER_REG_14__SCAN_IN) | (~new_n2653_ & ~P2_PHYADDRPOINTER_REG_14__SCAN_IN));
  assign new_n2653_ = P2_PHYADDRPOINTER_REG_13__SCAN_IN & new_n2020_ & P2_PHYADDRPOINTER_REG_10__SCAN_IN & new_n2019_ & P2_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign new_n2654_ = ~new_n2655_ & new_n4433_ & new_n4431_ & new_n2660_ & new_n2676_ & ~new_n4451_ & new_n2714_ & new_n4425_;
  assign new_n2655_ = (~new_n2596_ | (~new_n2656_ ^ (~new_n2561_ & (~new_n2521_ | ~new_n2560_)))) & new_n2657_ & (~new_n2564_ | ~new_n2659_);
  assign new_n2656_ = new_n2558_ ^ ~P1_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign new_n2657_ = (~P1_INSTADDRPOINTER_REG_23__SCAN_IN | (~new_n2574_ & (~new_n2586_ | (P1_INSTADDRPOINTER_REG_23__SCAN_IN & new_n2577_ & P1_INSTADDRPOINTER_REG_0__SCAN_IN)))) & new_n2658_ & (~new_n2577_ | ~P1_INSTADDRPOINTER_REG_0__SCAN_IN | ~new_n2586_ | (P1_INSTADDRPOINTER_REG_23__SCAN_IN & new_n2577_ & P1_INSTADDRPOINTER_REG_0__SCAN_IN)) & (~new_n2588_ | (~new_n2591_ & ~P1_INSTADDRPOINTER_REG_23__SCAN_IN) | (new_n2591_ & P1_INSTADDRPOINTER_REG_23__SCAN_IN));
  assign new_n2658_ = (~new_n2589_ | ~P1_REIP_REG_23__SCAN_IN) & ((~new_n2577_ & ~P1_INSTADDRPOINTER_REG_23__SCAN_IN) | ~new_n2584_ | (new_n2577_ & P1_INSTADDRPOINTER_REG_23__SCAN_IN));
  assign new_n2659_ = new_n2475_ ^ (new_n2472_ & ~new_n2474_ & new_n2453_ & new_n2473_);
  assign new_n2660_ = new_n2661_ & ((P2_INSTADDRPOINTER_REG_17__SCAN_IN & P2_INSTADDRPOINTER_REG_15__SCAN_IN & P2_INSTADDRPOINTER_REG_16__SCAN_IN & new_n1959_ & new_n1973_) | ~new_n2028_ | (~P2_INSTADDRPOINTER_REG_17__SCAN_IN & (~P2_INSTADDRPOINTER_REG_15__SCAN_IN | ~P2_INSTADDRPOINTER_REG_16__SCAN_IN | ~new_n1959_ | ~new_n1973_)));
  assign new_n2661_ = ~new_n2664_ & (((new_n2662_ | ~new_n2672_) & new_n2596_ & (~new_n2662_ | new_n2672_)) | ~new_n2675_ | new_n2673_ | ~new_n2674_);
  assign new_n2662_ = ~new_n2663_ & (new_n2549_ | (~new_n2523_ & (~new_n2548_ | (new_n2546_ & (new_n2524_ | new_n2530_)))));
  assign new_n2663_ = P1_INSTADDRPOINTER_REG_12__SCAN_IN & new_n2479_ & (~new_n2047_ | new_n2244_) & (new_n2047_ | ~new_n2244_);
  assign new_n2664_ = new_n2665_ & (~new_n2671_ | (~new_n1752_ & ~new_n1746_ & new_n1744_ & ~new_n1745_)) & (new_n2671_ | new_n1752_ | new_n1746_ | ~new_n1744_ | new_n1745_);
  assign new_n2665_ = new_n2669_ & new_n2666_ & P2_STATE2_REG_2__SCAN_IN & new_n2670_ & ~new_n1790_ & ~P2_STATEBS16_REG_SCAN_IN;
  assign new_n2666_ = new_n1791_ & ((~new_n2668_ & new_n1788_) | (new_n2667_ & ~new_n1762_ & (new_n1768_ | ~new_n1781_)));
  assign new_n2667_ = new_n1786_ & ~new_n1322_;
  assign new_n2668_ = (~new_n1786_ | ~new_n1322_) & (~new_n1787_ | new_n1370_);
  assign new_n2669_ = new_n1322_ & ~new_n1370_;
  assign new_n2670_ = ~new_n1378_ & ~P2_STATE_REG_0__SCAN_IN;
  assign new_n2671_ = (new_n1545_ | ~P2_INSTADDRPOINTER_REG_31__SCAN_IN) & (~new_n1542_ | ~P2_REIP_REG_31__SCAN_IN) & (~new_n1544_ | ~P2_EAX_REG_31__SCAN_IN);
  assign new_n2672_ = ~P1_INSTADDRPOINTER_REG_13__SCAN_IN ^ (~new_n2479_ | ((~new_n2227_ ^ ~new_n2163_) & new_n2047_ & (new_n2232_ ^ new_n2163_)) | ((~new_n2227_ | new_n2163_) & (new_n2227_ | ~new_n2163_) & (~new_n2047_ | (~new_n2232_ ^ new_n2163_))));
  assign new_n2673_ = new_n2588_ & (~P1_INSTADDRPOINTER_REG_13__SCAN_IN | ~new_n2594_ | ~P1_INSTADDRPOINTER_REG_8__SCAN_IN | ~P1_INSTADDRPOINTER_REG_10__SCAN_IN | ~P1_INSTADDRPOINTER_REG_9__SCAN_IN | ~P1_INSTADDRPOINTER_REG_12__SCAN_IN | ~P1_INSTADDRPOINTER_REG_11__SCAN_IN) & (P1_INSTADDRPOINTER_REG_13__SCAN_IN | (new_n2594_ & P1_INSTADDRPOINTER_REG_8__SCAN_IN & P1_INSTADDRPOINTER_REG_10__SCAN_IN & P1_INSTADDRPOINTER_REG_9__SCAN_IN & P1_INSTADDRPOINTER_REG_12__SCAN_IN & P1_INSTADDRPOINTER_REG_11__SCAN_IN));
  assign new_n2674_ = (~new_n2574_ | ~P1_INSTADDRPOINTER_REG_13__SCAN_IN) & (~new_n2564_ | (new_n2638_ & new_n2468_) | (~new_n2638_ & ~new_n2468_));
  assign new_n2675_ = (~new_n2589_ | ~P1_REIP_REG_13__SCAN_IN) & (~new_n2584_ | (~new_n2580_ & ~P1_INSTADDRPOINTER_REG_13__SCAN_IN) | (new_n2580_ & P1_INSTADDRPOINTER_REG_13__SCAN_IN)) & (~new_n2586_ | (~P1_INSTADDRPOINTER_REG_13__SCAN_IN & (~new_n2580_ | ~P1_INSTADDRPOINTER_REG_0__SCAN_IN)) | (P1_INSTADDRPOINTER_REG_0__SCAN_IN & new_n2580_ & P1_INSTADDRPOINTER_REG_13__SCAN_IN));
  assign new_n2676_ = new_n2694_ & ~new_n2677_ & ~new_n2679_ & ~new_n2681_ & ~new_n2703_ & ~new_n2688_ & (new_n2685_ | ~new_n2704_);
  assign new_n2677_ = new_n1751_ & new_n2678_;
  assign new_n2678_ = new_n1759_ & new_n1335_;
  assign new_n2679_ = (new_n2680_ | new_n2549_ | new_n2663_) & new_n2604_ & (~new_n2680_ | (~new_n2549_ & ~new_n2663_));
  assign new_n2680_ = ~new_n2523_ & (~new_n2548_ | (new_n2546_ & (new_n2524_ | new_n2530_)));
  assign new_n2681_ = (~new_n2683_ | new_n1335_ | (~new_n1707_ ^ (new_n1510_ & new_n1309_ & ~new_n1520_))) & (new_n2683_ | ~P2_EBX_REG_23__SCAN_IN) & (~new_n2682_ | ~new_n2683_ | ~new_n1335_);
  assign new_n2682_ = ~new_n2001_ ^ (new_n1976_ & ~new_n2000_);
  assign new_n2683_ = new_n1791_ & ((new_n1760_ & new_n1764_) | (new_n2684_ & (new_n1762_ | (~new_n1768_ & new_n1781_))));
  assign new_n2684_ = new_n1764_ & new_n1367_ & new_n1784_ & ~new_n1345_ & ~new_n1335_ & ~new_n1350_;
  assign new_n2685_ = (((new_n1960_ | P2_INSTADDRPOINTER_REG_6__SCAN_IN) & (new_n1961_ | (new_n1960_ & P2_INSTADDRPOINTER_REG_6__SCAN_IN))) | (new_n1799_ & P2_INSTADDRPOINTER_REG_7__SCAN_IN) | (~new_n1799_ & ~P2_INSTADDRPOINTER_REG_7__SCAN_IN)) & ~new_n2686_ & ~new_n2687_ & ((~new_n1960_ & ~P2_INSTADDRPOINTER_REG_6__SCAN_IN) | (~new_n1961_ & (~new_n1960_ | ~P2_INSTADDRPOINTER_REG_6__SCAN_IN)) | (new_n1799_ ^ P2_INSTADDRPOINTER_REG_7__SCAN_IN));
  assign new_n2686_ = ((new_n1963_ & P2_INSTADDRPOINTER_REG_4__SCAN_IN) | ((new_n1963_ | P2_INSTADDRPOINTER_REG_4__SCAN_IN) & ((new_n1964_ & P2_INSTADDRPOINTER_REG_3__SCAN_IN) | (new_n1965_ & (new_n1964_ | P2_INSTADDRPOINTER_REG_3__SCAN_IN))))) ^ (~new_n1962_ ^ ~P2_INSTADDRPOINTER_REG_5__SCAN_IN);
  assign new_n2687_ = ((new_n1968_ & P2_INSTADDRPOINTER_REG_1__SCAN_IN) | (new_n1966_ & (~new_n1587_ | ~new_n1322_ | ~new_n1580_) & (new_n1968_ | P2_INSTADDRPOINTER_REG_1__SCAN_IN))) ^ (P2_INSTADDRPOINTER_REG_2__SCAN_IN ^ (new_n1966_ ^ ~new_n1967_));
  assign new_n2688_ = (new_n2693_ | ~new_n2689_ | new_n2692_) & (new_n2690_ | new_n2691_) & (~new_n2693_ | (new_n2689_ & ~new_n2692_));
  assign new_n2689_ = ~new_n2027_ & new_n1975_ & new_n2023_;
  assign new_n2690_ = new_n2683_ & new_n1335_;
  assign new_n2691_ = ~new_n1790_ & ~P2_STATEBS16_REG_SCAN_IN & new_n1764_ & new_n2666_ & P2_STATE2_REG_2__SCAN_IN;
  assign new_n2692_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_30__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_30__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_30__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_30__SCAN_IN);
  assign new_n2693_ = (new_n1373_ | ~P2_INSTADDRPOINTER_REG_31__SCAN_IN) & (~new_n1380_ | ~P2_REIP_REG_31__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_31__SCAN_IN) & (~new_n1381_ | ~P2_EBX_REG_31__SCAN_IN);
  assign new_n2694_ = (~new_n2696_ | (new_n2649_ & (new_n2695_ | new_n2700_ | new_n2701_) & (~new_n2695_ | (~new_n2700_ & ~new_n2701_)))) & (~new_n2702_ | (new_n2503_ & (new_n2695_ | new_n2700_ | new_n2701_) & (~new_n2695_ | (~new_n2700_ & ~new_n2701_))));
  assign new_n2695_ = ~new_n2046_ & (new_n2242_ | (~new_n2243_ & (new_n2248_ | (~new_n2249_ & new_n2304_))));
  assign new_n2696_ = new_n2697_ & (~new_n2639_ | (P1_REIP_REG_14__SCAN_IN & new_n2646_ & P1_REIP_REG_13__SCAN_IN & P1_REIP_REG_12__SCAN_IN) | (~P1_REIP_REG_14__SCAN_IN & (~new_n2646_ | ~P1_REIP_REG_13__SCAN_IN | ~P1_REIP_REG_12__SCAN_IN)));
  assign new_n2697_ = (~new_n2643_ | (P1_PHYADDRPOINTER_REG_14__SCAN_IN & new_n2240_ & P1_PHYADDRPOINTER_REG_13__SCAN_IN) | (~P1_PHYADDRPOINTER_REG_14__SCAN_IN & (~new_n2240_ | ~P1_PHYADDRPOINTER_REG_13__SCAN_IN))) & new_n2698_ & (new_n2640_ | ~P1_EBX_REG_14__SCAN_IN);
  assign new_n2698_ = (~new_n2629_ | ~new_n2699_) & ~new_n2636_ & (~new_n2630_ | ~P1_REIP_REG_14__SCAN_IN) & (~P1_PHYADDRPOINTER_REG_14__SCAN_IN | new_n2630_ | ~P1_STATE2_REG_3__SCAN_IN);
  assign new_n2699_ = (new_n2638_ & new_n2468_) ^ (~new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_14__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_14__SCAN_IN)));
  assign new_n2700_ = new_n2322_ & (~new_n2237_ | (new_n2309_ & (new_n2311_ ^ new_n2163_)) | (~new_n2309_ & (new_n2311_ | ~new_n2163_) & (~new_n2311_ | new_n2163_)));
  assign new_n2701_ = ~new_n2322_ & new_n2237_ & (~new_n2309_ | (~new_n2311_ ^ new_n2163_)) & (new_n2309_ | (~new_n2311_ & new_n2163_) | (new_n2311_ & ~new_n2163_));
  assign new_n2702_ = (new_n2476_ | ~P1_EBX_REG_14__SCAN_IN) & (~new_n2699_ | ~new_n2476_ | ~new_n2053_);
  assign new_n2703_ = new_n2665_ & ((new_n1629_ ^ (new_n1628_ | new_n1627_ | ~new_n1528_ | new_n1626_)) | (new_n1528_ ^ ~new_n1626_));
  assign new_n2704_ = new_n2705_ & new_n2669_;
  assign new_n2705_ = new_n2706_ & new_n2708_;
  assign new_n2706_ = new_n1791_ & ((new_n2712_ & (new_n1762_ | (~new_n1768_ & new_n1781_))) | new_n2707_ | ~new_n2710_ | (new_n2713_ & ~new_n1762_ & (new_n1768_ | ~new_n1781_)));
  assign new_n2707_ = new_n2708_ & (new_n2709_ | (new_n2669_ & new_n2009_ & (~new_n1875_ | ~new_n1782_ | ~new_n2007_ | new_n2008_)));
  assign new_n2708_ = new_n1356_ & new_n1367_ & ~new_n1317_ & ~new_n1330_ & new_n1350_;
  assign new_n2709_ = ~new_n1322_ & new_n2011_;
  assign new_n2710_ = (~new_n1788_ | new_n1790_ | (new_n1322_ & new_n1367_) | (~new_n1787_ & ~new_n1322_)) & new_n2711_ & (~new_n1787_ | ~new_n1788_ | ~new_n2670_ | new_n1790_);
  assign new_n2711_ = ((~new_n1335_ & ~new_n1317_ & ~new_n1330_ & new_n1350_ & new_n1370_ & new_n1345_ & ~new_n1367_) | ((~new_n1370_ | (new_n1322_ & ~new_n1350_)) & (new_n1350_ | (~new_n1330_ & new_n1317_)) & ~new_n1335_ & ~new_n1345_ & new_n1367_)) & ((~new_n1330_ ^ new_n1317_) | (~new_n1330_ & ~new_n1350_)) & (~new_n1322_ | new_n1370_ | (~new_n1335_ & (new_n1330_ | ~new_n1317_) & (~new_n1330_ | new_n1317_)));
  assign new_n2712_ = ~new_n1370_ & ~new_n1350_;
  assign new_n2713_ = new_n1367_ ? (new_n1322_ & ~new_n1350_) : (~new_n1322_ & new_n2670_ & ~new_n1790_);
  assign new_n2714_ = ~new_n2715_ & new_n4414_ & new_n2716_ & new_n4354_ & ~new_n4421_ & new_n4351_ & new_n2758_ & new_n2771_;
  assign new_n2715_ = new_n2683_ & ~new_n1335_ & (new_n1704_ | ~new_n1509_ | (~new_n1703_ & (~new_n1510_ | ~new_n1309_ | new_n1520_))) & (~new_n1704_ | (new_n1509_ & (new_n1703_ | (new_n1510_ & new_n1309_ & ~new_n1520_))));
  assign new_n2716_ = (new_n2718_ | ~new_n2720_) & ~new_n2719_ & ((new_n2717_ & (new_n1650_ | new_n1686_) & (~new_n1650_ | ~new_n1686_)) | ~new_n1758_ | (~new_n2717_ & (new_n1650_ ^ ~new_n1686_)));
  assign new_n2717_ = ~new_n1652_ & (~new_n1685_ | (~new_n1655_ & new_n1682_));
  assign new_n2718_ = new_n2665_ & (new_n1628_ | new_n1627_ | ~new_n1528_ | new_n1626_) & (~new_n1628_ | (~new_n1627_ & new_n1528_ & ~new_n1626_));
  assign new_n2719_ = (new_n2243_ | new_n2248_ | (~new_n2249_ & new_n2304_)) & (new_n2602_ | new_n2649_) & ((~new_n2243_ & ~new_n2248_) | new_n2249_ | ~new_n2304_);
  assign new_n2720_ = (~new_n2691_ | (~new_n2002_ & ~new_n2001_ & new_n1976_ & ~new_n2000_) | (new_n2002_ & (new_n2001_ | ~new_n1976_ | new_n2000_))) & new_n2721_ & (~new_n1946_ | ~new_n2757_);
  assign new_n2721_ = (~new_n2726_ | ~new_n2729_) & new_n2722_ & (~new_n2756_ | (new_n2017_ & P2_PHYADDRPOINTER_REG_24__SCAN_IN) | (~new_n2017_ & ~P2_PHYADDRPOINTER_REG_24__SCAN_IN));
  assign new_n2722_ = (new_n2723_ | ~P2_EBX_REG_24__SCAN_IN) & (~new_n2724_ | ~P2_REIP_REG_24__SCAN_IN) & (~P2_PHYADDRPOINTER_REG_24__SCAN_IN | new_n2724_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n2723_ = (P2_EBX_REG_31__SCAN_IN | (~new_n1790_ & ~P2_STATEBS16_REG_SCAN_IN) | new_n1322_ | new_n1370_ | ~new_n2666_ | ~P2_STATE2_REG_2__SCAN_IN) & (~new_n1322_ | new_n1370_ | ~new_n2666_ | ~P2_STATE2_REG_2__SCAN_IN | (new_n2670_ & ~new_n1790_ & ~P2_STATEBS16_REG_SCAN_IN));
  assign new_n2724_ = new_n2725_ & (~new_n1791_ | ((new_n2668_ | ~new_n1788_) & (~new_n2667_ | new_n1762_ | (~new_n1768_ & new_n1781_))));
  assign new_n2725_ = (~P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_1__SCAN_IN | P2_STATE2_REG_2__SCAN_IN | ~P2_STATE2_REG_0__SCAN_IN) & (P2_STATE2_REG_2__SCAN_IN | P2_STATE2_REG_1__SCAN_IN | P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_0__SCAN_IN) & (~P2_STATE2_REG_1__SCAN_IN | P2_STATEBS16_REG_SCAN_IN | P2_STATE2_REG_2__SCAN_IN | P2_STATE2_REG_0__SCAN_IN);
  assign new_n2726_ = ~new_n2727_ & ~new_n2724_ & P2_STATE2_REG_1__SCAN_IN;
  assign new_n2727_ = P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_31__SCAN_IN : (~new_n2728_ ^ P2_PHYADDRPOINTER_REG_31__SCAN_IN);
  assign new_n2728_ = P2_PHYADDRPOINTER_REG_30__SCAN_IN & P2_PHYADDRPOINTER_REG_29__SCAN_IN & P2_PHYADDRPOINTER_REG_28__SCAN_IN & P2_PHYADDRPOINTER_REG_26__SCAN_IN & P2_PHYADDRPOINTER_REG_27__SCAN_IN & P2_PHYADDRPOINTER_REG_25__SCAN_IN & new_n2017_ & P2_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign new_n2729_ = (P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_24__SCAN_IN : (~P2_PHYADDRPOINTER_REG_24__SCAN_IN ^ (new_n2730_ & P2_PHYADDRPOINTER_REG_23__SCAN_IN))) ^ (new_n2733_ & new_n2755_ & (~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN) & (P2_STATE2_REG_0__SCAN_IN | (~new_n2730_ & ~P2_PHYADDRPOINTER_REG_23__SCAN_IN) | (new_n2730_ & P2_PHYADDRPOINTER_REG_23__SCAN_IN)));
  assign new_n2730_ = P2_PHYADDRPOINTER_REG_22__SCAN_IN & new_n2731_ & P2_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign new_n2731_ = P2_PHYADDRPOINTER_REG_20__SCAN_IN & P2_PHYADDRPOINTER_REG_19__SCAN_IN & new_n2732_ & P2_PHYADDRPOINTER_REG_18__SCAN_IN;
  assign new_n2732_ = new_n2018_ & P2_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign new_n2733_ = new_n2754_ & new_n2734_ & new_n2753_ & new_n2735_ & new_n2736_ & new_n2751_;
  assign new_n2734_ = P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_20__SCAN_IN : (~P2_PHYADDRPOINTER_REG_20__SCAN_IN ^ (P2_PHYADDRPOINTER_REG_19__SCAN_IN & new_n2732_ & P2_PHYADDRPOINTER_REG_18__SCAN_IN));
  assign new_n2735_ = P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_18__SCAN_IN : (~new_n2732_ ^ P2_PHYADDRPOINTER_REG_18__SCAN_IN);
  assign new_n2736_ = ~new_n2737_ & ~new_n2750_ & new_n2746_ & ~new_n2744_ & ~new_n2749_ & new_n2747_ & new_n2738_ & ~new_n2748_;
  assign new_n2737_ = ~P2_STATE2_REG_0__SCAN_IN & (~P2_PHYADDRPOINTER_REG_15__SCAN_IN | ~new_n2653_ | ~P2_PHYADDRPOINTER_REG_14__SCAN_IN) & (P2_PHYADDRPOINTER_REG_15__SCAN_IN | (new_n2653_ & P2_PHYADDRPOINTER_REG_14__SCAN_IN));
  assign new_n2738_ = ~new_n2741_ & (~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_6__SCAN_IN) & (P2_STATE2_REG_0__SCAN_IN | (P2_PHYADDRPOINTER_REG_6__SCAN_IN & new_n2743_ & P2_PHYADDRPOINTER_REG_5__SCAN_IN) | (~P2_PHYADDRPOINTER_REG_6__SCAN_IN & (~new_n2743_ | ~P2_PHYADDRPOINTER_REG_5__SCAN_IN))) & new_n2739_ & (~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_5__SCAN_IN) & (P2_STATE2_REG_0__SCAN_IN | (new_n2743_ & P2_PHYADDRPOINTER_REG_5__SCAN_IN) | (~new_n2743_ & ~P2_PHYADDRPOINTER_REG_5__SCAN_IN));
  assign new_n2739_ = (~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_4__SCAN_IN) & (P2_STATE2_REG_0__SCAN_IN | (P2_PHYADDRPOINTER_REG_4__SCAN_IN & P2_PHYADDRPOINTER_REG_3__SCAN_IN & P2_PHYADDRPOINTER_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_2__SCAN_IN) | (~P2_PHYADDRPOINTER_REG_4__SCAN_IN & (~P2_PHYADDRPOINTER_REG_3__SCAN_IN | ~P2_PHYADDRPOINTER_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_2__SCAN_IN))) & new_n2740_ & (~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_3__SCAN_IN) & ((~P2_PHYADDRPOINTER_REG_3__SCAN_IN & (~P2_PHYADDRPOINTER_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_2__SCAN_IN)) | P2_STATE2_REG_0__SCAN_IN | (P2_PHYADDRPOINTER_REG_3__SCAN_IN & P2_PHYADDRPOINTER_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_2__SCAN_IN));
  assign new_n2740_ = (P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_0__SCAN_IN : ~P2_PHYADDRPOINTER_REG_0__SCAN_IN) & (P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_1__SCAN_IN : P2_PHYADDRPOINTER_REG_1__SCAN_IN) & (~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_2__SCAN_IN) & (P2_STATE2_REG_0__SCAN_IN | (~P2_PHYADDRPOINTER_REG_1__SCAN_IN & ~P2_PHYADDRPOINTER_REG_2__SCAN_IN) | (P2_PHYADDRPOINTER_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_2__SCAN_IN));
  assign new_n2741_ = (new_n2742_ | P2_STATE2_REG_0__SCAN_IN) & (P2_INSTADDRPOINTER_REG_8__SCAN_IN | P2_INSTADDRPOINTER_REG_9__SCAN_IN | ~P2_STATE2_REG_0__SCAN_IN | P2_INSTADDRPOINTER_REG_7__SCAN_IN);
  assign new_n2742_ = (~P2_PHYADDRPOINTER_REG_8__SCAN_IN | ~P2_PHYADDRPOINTER_REG_7__SCAN_IN | ~P2_PHYADDRPOINTER_REG_6__SCAN_IN | ~P2_PHYADDRPOINTER_REG_5__SCAN_IN | ~P2_PHYADDRPOINTER_REG_4__SCAN_IN | ~P2_PHYADDRPOINTER_REG_3__SCAN_IN | ~P2_PHYADDRPOINTER_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_2__SCAN_IN) & (P2_PHYADDRPOINTER_REG_7__SCAN_IN | P2_PHYADDRPOINTER_REG_8__SCAN_IN | (P2_PHYADDRPOINTER_REG_6__SCAN_IN & P2_PHYADDRPOINTER_REG_5__SCAN_IN & P2_PHYADDRPOINTER_REG_4__SCAN_IN & P2_PHYADDRPOINTER_REG_3__SCAN_IN & P2_PHYADDRPOINTER_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_2__SCAN_IN));
  assign new_n2743_ = P2_PHYADDRPOINTER_REG_4__SCAN_IN & P2_PHYADDRPOINTER_REG_3__SCAN_IN & P2_PHYADDRPOINTER_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign new_n2744_ = P2_STATE2_REG_0__SCAN_IN ? P2_INSTADDRPOINTER_REG_13__SCAN_IN : (new_n2745_ ^ P2_PHYADDRPOINTER_REG_13__SCAN_IN);
  assign new_n2745_ = new_n2020_ & P2_PHYADDRPOINTER_REG_10__SCAN_IN & new_n2019_ & P2_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign new_n2746_ = P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_14__SCAN_IN : (~new_n2653_ ^ P2_PHYADDRPOINTER_REG_14__SCAN_IN);
  assign new_n2747_ = P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_10__SCAN_IN : (P2_PHYADDRPOINTER_REG_10__SCAN_IN ^ (~new_n2019_ | ~P2_PHYADDRPOINTER_REG_9__SCAN_IN));
  assign new_n2748_ = (new_n2019_ | P2_PHYADDRPOINTER_REG_9__SCAN_IN) & ~P2_STATE2_REG_0__SCAN_IN & (~new_n2019_ | ~P2_PHYADDRPOINTER_REG_9__SCAN_IN);
  assign new_n2749_ = (P2_INSTADDRPOINTER_REG_12__SCAN_IN | ~P2_STATE2_REG_0__SCAN_IN | P2_INSTADDRPOINTER_REG_11__SCAN_IN) & (P2_STATE2_REG_0__SCAN_IN | ((P2_PHYADDRPOINTER_REG_10__SCAN_IN & new_n2019_ & P2_PHYADDRPOINTER_REG_9__SCAN_IN) ? (~P2_PHYADDRPOINTER_REG_11__SCAN_IN | ~P2_PHYADDRPOINTER_REG_12__SCAN_IN) : (P2_PHYADDRPOINTER_REG_11__SCAN_IN | P2_PHYADDRPOINTER_REG_12__SCAN_IN)));
  assign new_n2750_ = P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign new_n2751_ = (~P2_STATE2_REG_0__SCAN_IN | (~P2_INSTADDRPOINTER_REG_16__SCAN_IN & ~P2_INSTADDRPOINTER_REG_17__SCAN_IN)) & ((P2_PHYADDRPOINTER_REG_17__SCAN_IN & new_n2752_ & P2_PHYADDRPOINTER_REG_16__SCAN_IN) | P2_STATE2_REG_0__SCAN_IN | (~new_n2752_ & ~P2_PHYADDRPOINTER_REG_16__SCAN_IN & ~P2_PHYADDRPOINTER_REG_17__SCAN_IN));
  assign new_n2752_ = P2_PHYADDRPOINTER_REG_15__SCAN_IN & new_n2653_ & P2_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign new_n2753_ = (~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_19__SCAN_IN) & ((~P2_PHYADDRPOINTER_REG_19__SCAN_IN & (~new_n2732_ | ~P2_PHYADDRPOINTER_REG_18__SCAN_IN)) | P2_STATE2_REG_0__SCAN_IN | (P2_PHYADDRPOINTER_REG_19__SCAN_IN & new_n2732_ & P2_PHYADDRPOINTER_REG_18__SCAN_IN));
  assign new_n2754_ = P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_21__SCAN_IN : (~P2_PHYADDRPOINTER_REG_21__SCAN_IN ^ (P2_PHYADDRPOINTER_REG_20__SCAN_IN & P2_PHYADDRPOINTER_REG_19__SCAN_IN & new_n2732_ & P2_PHYADDRPOINTER_REG_18__SCAN_IN));
  assign new_n2755_ = P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_22__SCAN_IN : (P2_PHYADDRPOINTER_REG_22__SCAN_IN ^ (~new_n2731_ | ~P2_PHYADDRPOINTER_REG_21__SCAN_IN));
  assign new_n2756_ = new_n2727_ & ~new_n2724_ & P2_STATE2_REG_1__SCAN_IN;
  assign new_n2757_ = P2_EBX_REG_31__SCAN_IN & (new_n1790_ | P2_STATEBS16_REG_SCAN_IN) & new_n1764_ & new_n2666_ & P2_STATE2_REG_2__SCAN_IN;
  assign new_n2758_ = ~new_n2759_ & ~new_n2766_ & (~new_n2691_ | (~new_n2003_ & ~new_n2002_ & ~new_n2001_ & new_n1976_ & ~new_n2000_) | (new_n2003_ & (new_n2002_ | new_n2001_ | ~new_n1976_ | new_n2000_)));
  assign new_n2759_ = (~new_n1639_ | ~new_n2665_) & new_n2760_ & ((new_n1999_ & (new_n1998_ | ~new_n2765_ | new_n1997_)) | ~new_n2691_ | (~new_n1999_ & ~new_n1998_ & new_n2765_ & ~new_n1997_));
  assign new_n2760_ = new_n2761_ & (~new_n2757_ | (new_n1330_ & P2_EBX_REG_21__SCAN_IN & (~new_n1942_ | (new_n1330_ & P2_EBX_REG_19__SCAN_IN) | new_n1907_ | (new_n1330_ & P2_EBX_REG_20__SCAN_IN))) | new_n1907_ | ((~new_n1330_ | ~P2_EBX_REG_21__SCAN_IN) & new_n1942_ & (~new_n1330_ | ~P2_EBX_REG_19__SCAN_IN) & ~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_20__SCAN_IN)));
  assign new_n2761_ = (~new_n2726_ | (new_n2763_ & (~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_21__SCAN_IN) & (P2_STATE2_REG_0__SCAN_IN | (new_n2731_ & P2_PHYADDRPOINTER_REG_21__SCAN_IN) | (~new_n2731_ & ~P2_PHYADDRPOINTER_REG_21__SCAN_IN))) | (~new_n2763_ & (P2_STATE2_REG_0__SCAN_IN ? P2_INSTADDRPOINTER_REG_21__SCAN_IN : (new_n2731_ ^ P2_PHYADDRPOINTER_REG_21__SCAN_IN)))) & new_n2762_ & (~new_n2756_ | (new_n2731_ & P2_PHYADDRPOINTER_REG_21__SCAN_IN) | (~new_n2731_ & ~P2_PHYADDRPOINTER_REG_21__SCAN_IN));
  assign new_n2762_ = (new_n2723_ | ~P2_EBX_REG_21__SCAN_IN) & (~new_n2724_ | ~P2_REIP_REG_21__SCAN_IN) & (~P2_PHYADDRPOINTER_REG_21__SCAN_IN | new_n2724_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n2763_ = new_n2734_ & new_n2764_ & new_n2753_;
  assign new_n2764_ = new_n2735_ & new_n2736_ & new_n2751_;
  assign new_n2765_ = ~new_n1996_ & ~new_n1995_ & ~new_n1994_ & new_n1977_ & ~new_n1993_;
  assign new_n2766_ = ~new_n2767_ & new_n2768_ & ((~P1_INSTADDRPOINTER_REG_6__SCAN_IN & (~new_n2582_ | (~new_n2584_ & ~P1_INSTADDRPOINTER_REG_0__SCAN_IN))) | (~new_n2584_ & ~new_n2586_) | (new_n2582_ & P1_INSTADDRPOINTER_REG_6__SCAN_IN & (~new_n2586_ | P1_INSTADDRPOINTER_REG_0__SCAN_IN)));
  assign new_n2767_ = new_n2596_ & ((~new_n2533_ & P1_INSTADDRPOINTER_REG_6__SCAN_IN) | (new_n2533_ & ~P1_INSTADDRPOINTER_REG_6__SCAN_IN) | ((new_n2534_ | ~P1_INSTADDRPOINTER_REG_5__SCAN_IN) & (new_n2535_ | (new_n2534_ & ~P1_INSTADDRPOINTER_REG_5__SCAN_IN)))) & ((~new_n2533_ ^ P1_INSTADDRPOINTER_REG_6__SCAN_IN) | (~new_n2534_ & P1_INSTADDRPOINTER_REG_5__SCAN_IN) | (~new_n2535_ & (~new_n2534_ | P1_INSTADDRPOINTER_REG_5__SCAN_IN)));
  assign new_n2768_ = (~P1_REIP_REG_6__SCAN_IN | new_n2574_ | P1_STATE2_REG_2__SCAN_IN) & (~new_n2588_ | (new_n2595_ & P1_INSTADDRPOINTER_REG_6__SCAN_IN) | (~new_n2595_ & ~P1_INSTADDRPOINTER_REG_6__SCAN_IN)) & (~new_n2564_ | ~new_n2769_) & (~new_n2574_ | ~P1_INSTADDRPOINTER_REG_6__SCAN_IN);
  assign new_n2769_ = (~new_n2770_ | new_n2461_) ^ (new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_6__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_6__SCAN_IN)));
  assign new_n2770_ = ~new_n2458_ & ~new_n2459_ & ~new_n2460_;
  assign new_n2771_ = new_n4344_ & new_n2772_ & new_n4237_ & new_n4186_ & new_n2959_ & new_n4128_ & new_n3110_ & new_n3225_;
  assign new_n2772_ = new_n2774_ & ~new_n2951_ & (((~new_n2773_ | new_n1907_ | (new_n1330_ & P2_EBX_REG_30__SCAN_IN)) & (new_n1907_ | (new_n1330_ & P2_EBX_REG_31__SCAN_IN))) | ~new_n2757_ | (~new_n1330_ & new_n2773_ & ~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_30__SCAN_IN)));
  assign new_n2773_ = new_n2032_ & (~new_n1330_ | ~P2_EBX_REG_29__SCAN_IN);
  assign new_n2774_ = (~new_n1700_ | ~new_n2665_) & (~new_n2937_ | (new_n2775_ & ~new_n2929_));
  assign new_n2775_ = ((~P3_INSTADDRPOINTER_REG_25__SCAN_IN & (~P3_INSTADDRPOINTER_REG_24__SCAN_IN | ~new_n2863_ | ~P3_INSTADDRPOINTER_REG_23__SCAN_IN)) | ~new_n2928_ | (P3_INSTADDRPOINTER_REG_25__SCAN_IN & P3_INSTADDRPOINTER_REG_24__SCAN_IN & new_n2863_ & P3_INSTADDRPOINTER_REG_23__SCAN_IN)) & ((~P3_INSTADDRPOINTER_REG_25__SCAN_IN & (~P3_INSTADDRPOINTER_REG_24__SCAN_IN | ~new_n2911_ | ~P3_INSTADDRPOINTER_REG_23__SCAN_IN)) | ~new_n2926_ | (P3_INSTADDRPOINTER_REG_25__SCAN_IN & P3_INSTADDRPOINTER_REG_24__SCAN_IN & new_n2911_ & P3_INSTADDRPOINTER_REG_23__SCAN_IN)) & (~new_n2928_ | (new_n2863_ & P3_INSTADDRPOINTER_REG_23__SCAN_IN) | (~new_n2863_ & ~P3_INSTADDRPOINTER_REG_23__SCAN_IN)) & new_n2776_ & ((~new_n2911_ & ~P3_INSTADDRPOINTER_REG_23__SCAN_IN) | ~new_n2926_ | (new_n2911_ & P3_INSTADDRPOINTER_REG_23__SCAN_IN));
  assign new_n2776_ = ~new_n2855_ & ((~new_n2845_ & new_n2861_) | (P3_INSTADDRPOINTER_REG_25__SCAN_IN & new_n2851_ & P3_INSTADDRPOINTER_REG_0__SCAN_IN) | (~P3_INSTADDRPOINTER_REG_25__SCAN_IN & (~new_n2851_ | ~P3_INSTADDRPOINTER_REG_0__SCAN_IN))) & new_n2777_ & (new_n2862_ | (P3_INSTADDRPOINTER_REG_25__SCAN_IN & new_n2851_ & P3_INSTADDRPOINTER_REG_0__SCAN_IN) | (~P3_INSTADDRPOINTER_REG_25__SCAN_IN & (~new_n2851_ | ~P3_INSTADDRPOINTER_REG_0__SCAN_IN)));
  assign new_n2777_ = new_n2778_ & ~new_n2852_ & new_n2841_ & ((~new_n2839_ & ~new_n2840_) | (new_n2851_ & P3_INSTADDRPOINTER_REG_25__SCAN_IN) | (~new_n2851_ & ~P3_INSTADDRPOINTER_REG_25__SCAN_IN));
  assign new_n2778_ = ((~new_n2832_ & ~new_n2839_) | (new_n2779_ & P3_INSTADDRPOINTER_REG_23__SCAN_IN) | (~new_n2779_ & ~P3_INSTADDRPOINTER_REG_23__SCAN_IN)) & ((~new_n2788_ & ~new_n2840_) | (new_n2779_ & P3_INSTADDRPOINTER_REG_23__SCAN_IN) | (~new_n2779_ & ~P3_INSTADDRPOINTER_REG_23__SCAN_IN)) & ((~new_n2788_ & ~new_n2832_) | (P3_INSTADDRPOINTER_REG_25__SCAN_IN & P3_INSTADDRPOINTER_REG_24__SCAN_IN & new_n2779_ & P3_INSTADDRPOINTER_REG_23__SCAN_IN) | (~P3_INSTADDRPOINTER_REG_25__SCAN_IN & (~P3_INSTADDRPOINTER_REG_24__SCAN_IN | ~new_n2779_ | ~P3_INSTADDRPOINTER_REG_23__SCAN_IN)));
  assign new_n2779_ = P3_INSTADDRPOINTER_REG_22__SCAN_IN & new_n2780_ & new_n2786_;
  assign new_n2780_ = new_n2781_ & new_n2783_ & new_n2785_;
  assign new_n2781_ = new_n2782_ & P3_INSTADDRPOINTER_REG_15__SCAN_IN & P3_INSTADDRPOINTER_REG_17__SCAN_IN & P3_INSTADDRPOINTER_REG_16__SCAN_IN & P3_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign new_n2782_ = P3_INSTADDRPOINTER_REG_10__SCAN_IN & P3_INSTADDRPOINTER_REG_11__SCAN_IN & P3_INSTADDRPOINTER_REG_14__SCAN_IN & P3_INSTADDRPOINTER_REG_12__SCAN_IN & P3_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign new_n2783_ = new_n2784_ & P3_INSTADDRPOINTER_REG_3__SCAN_IN & P3_INSTADDRPOINTER_REG_4__SCAN_IN & P3_INSTADDRPOINTER_REG_7__SCAN_IN & P3_INSTADDRPOINTER_REG_5__SCAN_IN & P3_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign new_n2784_ = P3_INSTADDRPOINTER_REG_8__SCAN_IN & P3_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign new_n2785_ = P3_INSTADDRPOINTER_REG_1__SCAN_IN & P3_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign new_n2786_ = new_n2787_ & P3_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign new_n2787_ = P3_INSTADDRPOINTER_REG_19__SCAN_IN & P3_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign new_n2788_ = new_n2789_ & ~new_n2826_;
  assign new_n2789_ = new_n2802_ & new_n2809_ & new_n2815_ & new_n2821_ & ~new_n2790_ & new_n2796_;
  assign new_n2790_ = new_n2791_ & new_n2792_ & new_n2793_ & new_n2794_ & new_n2795_;
  assign new_n2791_ = (~P3_INSTQUEUE_REG_14__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_11__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2792_ = (~P3_INSTQUEUE_REG_7__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_15__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2793_ = (~P3_INSTQUEUE_REG_1__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2794_ = (~P3_INSTQUEUE_REG_10__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_0__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2795_ = (~P3_INSTQUEUE_REG_5__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_3__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2796_ = new_n2797_ & new_n2798_ & new_n2799_ & new_n2800_ & new_n2801_;
  assign new_n2797_ = (~P3_INSTQUEUE_REG_14__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_11__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2798_ = (~P3_INSTQUEUE_REG_7__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_15__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2799_ = (~P3_INSTQUEUE_REG_1__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2800_ = (~P3_INSTQUEUE_REG_10__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_0__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2801_ = (~P3_INSTQUEUE_REG_5__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_3__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2802_ = new_n2806_ & new_n2807_ & new_n2808_ & new_n2805_ & (~new_n2803_ | ~P3_INSTQUEUE_REG_7__1__SCAN_IN) & (~new_n2804_ | ~P3_INSTQUEUE_REG_15__1__SCAN_IN);
  assign new_n2803_ = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign new_n2804_ = P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign new_n2805_ = (~P3_INSTQUEUE_REG_14__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_11__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2806_ = (~P3_INSTQUEUE_REG_1__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2807_ = (~P3_INSTQUEUE_REG_10__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_0__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2808_ = (~P3_INSTQUEUE_REG_5__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_3__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2809_ = new_n2810_ & new_n2811_ & new_n2812_ & new_n2813_ & new_n2814_;
  assign new_n2810_ = (~P3_INSTQUEUE_REG_14__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_11__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2811_ = (~P3_INSTQUEUE_REG_7__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_15__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2812_ = (~P3_INSTQUEUE_REG_1__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2813_ = (~P3_INSTQUEUE_REG_10__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_0__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2814_ = (~P3_INSTQUEUE_REG_5__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_3__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2815_ = new_n2816_ & new_n2817_ & new_n2818_ & new_n2819_ & new_n2820_;
  assign new_n2816_ = (~P3_INSTQUEUE_REG_14__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_11__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2817_ = (~P3_INSTQUEUE_REG_7__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_15__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2818_ = (~P3_INSTQUEUE_REG_1__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2819_ = (~P3_INSTQUEUE_REG_10__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_0__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2820_ = (~P3_INSTQUEUE_REG_5__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_3__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2821_ = new_n2823_ & new_n2824_ & new_n2825_ & new_n2822_ & (~new_n2803_ | ~P3_INSTQUEUE_REG_7__3__SCAN_IN) & (~new_n2804_ | ~P3_INSTQUEUE_REG_15__3__SCAN_IN);
  assign new_n2822_ = (~P3_INSTQUEUE_REG_14__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_11__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2823_ = (~P3_INSTQUEUE_REG_1__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2824_ = (~P3_INSTQUEUE_REG_10__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_0__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2825_ = (~P3_INSTQUEUE_REG_5__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_3__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2826_ = new_n2827_ & new_n2828_ & new_n2829_ & new_n2830_ & new_n2831_;
  assign new_n2827_ = (~P3_INSTQUEUE_REG_14__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_11__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2828_ = (~P3_INSTQUEUE_REG_7__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_15__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2829_ = (~P3_INSTQUEUE_REG_1__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2830_ = (~P3_INSTQUEUE_REG_10__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_0__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2831_ = (~P3_INSTQUEUE_REG_5__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_3__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2832_ = new_n2802_ & new_n2833_ & ~new_n2790_ & ~new_n2796_ & ~new_n2826_ & new_n2821_ & new_n2809_ & ~new_n2815_;
  assign new_n2833_ = new_n2834_ & new_n2835_ & new_n2836_ & new_n2837_ & new_n2838_;
  assign new_n2834_ = (~P3_INSTQUEUE_REG_14__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_11__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2835_ = (~P3_INSTQUEUE_REG_7__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_15__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2836_ = (~P3_INSTQUEUE_REG_1__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2837_ = (~P3_INSTQUEUE_REG_10__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_0__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2838_ = (~P3_INSTQUEUE_REG_5__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_3__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2839_ = new_n2796_ & ~new_n2809_ & new_n2790_ & new_n2833_ & new_n2815_ & ~new_n2826_ & ~new_n2821_;
  assign new_n2840_ = ~new_n2826_ & new_n2821_ & new_n2833_ & ~new_n2790_ & ~new_n2796_ & ~new_n2815_ & ~new_n2802_ & new_n2809_;
  assign new_n2841_ = (~new_n2845_ | (new_n2842_ & P3_INSTADDRPOINTER_REG_23__SCAN_IN) | (~new_n2842_ & ~P3_INSTADDRPOINTER_REG_23__SCAN_IN)) & (~new_n2850_ | (~new_n2847_ & ~P3_INSTADDRPOINTER_REG_25__SCAN_IN) | (new_n2847_ & P3_INSTADDRPOINTER_REG_25__SCAN_IN));
  assign new_n2842_ = P3_INSTADDRPOINTER_REG_22__SCAN_IN & new_n2843_ & new_n2786_;
  assign new_n2843_ = new_n2781_ & new_n2783_ & new_n2844_;
  assign new_n2844_ = P3_INSTADDRPOINTER_REG_2__SCAN_IN & P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign new_n2845_ = new_n2846_ & new_n2809_;
  assign new_n2846_ = new_n2802_ & new_n2790_ & new_n2821_ & new_n2826_ & new_n2833_ & new_n2796_ & ~new_n2815_;
  assign new_n2847_ = P3_INSTADDRPOINTER_REG_24__SCAN_IN & P3_INSTADDRPOINTER_REG_23__SCAN_IN & P3_INSTADDRPOINTER_REG_22__SCAN_IN & new_n2848_ & new_n2786_;
  assign new_n2848_ = new_n2781_ & new_n2783_ & ~new_n2849_;
  assign new_n2849_ = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN & (~P3_INSTADDRPOINTER_REG_0__SCAN_IN | ~P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  assign new_n2850_ = (~new_n2802_ ^ new_n2809_) & ~new_n2826_ & ~new_n2821_ & new_n2790_ & ~new_n2796_ & new_n2815_ & ~new_n2833_;
  assign new_n2851_ = P3_INSTADDRPOINTER_REG_24__SCAN_IN & P3_INSTADDRPOINTER_REG_23__SCAN_IN & P3_INSTADDRPOINTER_REG_22__SCAN_IN & new_n2780_ & new_n2786_;
  assign new_n2852_ = (new_n2853_ | new_n2854_) & (~P3_INSTADDRPOINTER_REG_23__SCAN_IN | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN | ~new_n2848_ | ~new_n2786_) & (P3_INSTADDRPOINTER_REG_23__SCAN_IN | (P3_INSTADDRPOINTER_REG_22__SCAN_IN & new_n2848_ & new_n2786_));
  assign new_n2853_ = ~new_n2821_ & new_n2790_ & ~new_n2796_ & new_n2802_ & new_n2809_ & ~new_n2826_ & new_n2815_ & ~new_n2833_;
  assign new_n2854_ = ~new_n2802_ & ~new_n2809_ & ~new_n2826_ & ~new_n2821_ & new_n2790_ & ~new_n2796_ & new_n2815_ & ~new_n2833_;
  assign new_n2855_ = ~new_n2856_ & (new_n2779_ | P3_INSTADDRPOINTER_REG_23__SCAN_IN) & (P3_INSTADDRPOINTER_REG_0__SCAN_IN | P3_INSTADDRPOINTER_REG_23__SCAN_IN) & (~new_n2842_ | ~P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  assign new_n2856_ = new_n2857_ & ~new_n2858_ & ~new_n2859_ & new_n2860_ & (~new_n2846_ | new_n2809_);
  assign new_n2857_ = (~new_n2815_ | ((~new_n2802_ | new_n2809_ | (~new_n2821_ & (~new_n2790_ | new_n2796_) & ~new_n2826_ & (new_n2790_ | ~new_n2796_))) & (~new_n2809_ | ((~new_n2790_ | ~new_n2833_) & (~new_n2802_ | new_n2790_ | new_n2796_))) & ((new_n2796_ & new_n2826_) | new_n2802_ | (~new_n2826_ & ~new_n2821_)))) & (new_n2796_ | ~new_n2821_ | (new_n2809_ & (~new_n2802_ | ~new_n2826_))) & (new_n2796_ | new_n2802_ | ~new_n2790_ | ~new_n2833_) & (new_n2802_ | ~new_n2790_ | ~new_n2826_) & ((~new_n2790_ & ~new_n2796_) | new_n2802_ | ~new_n2809_) & (~new_n2796_ | new_n2821_ | (new_n2790_ & new_n2833_)) & (new_n2833_ | ((~new_n2802_ | new_n2809_) & ~new_n2826_ & (new_n2790_ | new_n2796_))) & (new_n2815_ | (new_n2821_ & (new_n2790_ ? new_n2826_ : ~new_n2796_))) & (new_n2802_ | new_n2809_ | ~new_n2826_ | ~new_n2833_ | ~new_n2815_ | ~new_n2821_ | new_n2790_ | ~new_n2796_);
  assign new_n2858_ = new_n2790_ & new_n2821_ & new_n2802_ & new_n2809_ & ~new_n2826_ & new_n2815_ & ~new_n2833_;
  assign new_n2859_ = new_n2826_ & new_n2821_ & new_n2833_ & ~new_n2790_ & ~new_n2796_ & ~new_n2815_ & ~new_n2802_ & new_n2809_;
  assign new_n2860_ = (new_n2802_ | ~new_n2809_ | ~new_n2833_ | new_n2790_ | new_n2796_ | ~new_n2815_ | new_n2826_ | new_n2821_) & (~new_n2826_ | ~new_n2833_ | ~new_n2802_ | ~new_n2809_ | ~new_n2815_ | ~new_n2821_ | new_n2790_ | ~new_n2796_);
  assign new_n2861_ = (~new_n2815_ | ((~new_n2802_ | new_n2809_ | (~new_n2821_ & (~new_n2790_ | new_n2796_) & ~new_n2826_ & (new_n2790_ | ~new_n2796_))) & (~new_n2809_ | ((~new_n2790_ | ~new_n2833_) & (~new_n2802_ | new_n2790_ | new_n2796_))) & ((new_n2796_ & new_n2826_) | new_n2802_ | (~new_n2826_ & ~new_n2821_)))) & (new_n2796_ | ~new_n2821_ | (new_n2809_ & (~new_n2802_ | ~new_n2826_))) & (new_n2796_ | new_n2802_ | ~new_n2790_ | ~new_n2833_) & (new_n2802_ | ~new_n2790_ | ~new_n2826_) & ((~new_n2790_ & ~new_n2796_) | new_n2802_ | ~new_n2809_) & (~new_n2796_ | new_n2821_ | (new_n2790_ & new_n2833_)) & (new_n2833_ | ((~new_n2802_ | new_n2809_) & ~new_n2826_ & (new_n2790_ | new_n2796_))) & (new_n2815_ | (new_n2821_ & (new_n2790_ ? new_n2826_ : ~new_n2796_)));
  assign new_n2862_ = ((new_n2802_ ^ new_n2809_) | ~new_n2826_ | ~new_n2833_ | ~new_n2815_ | ~new_n2821_ | new_n2790_ | ~new_n2796_) & (new_n2809_ | ~new_n2802_ | ~new_n2790_ | ~new_n2821_ | ~new_n2826_ | ~new_n2833_ | ~new_n2796_ | new_n2815_) & (new_n2802_ | ~new_n2809_ | ~new_n2833_ | new_n2790_ | new_n2796_ | ~new_n2815_ | new_n2826_ | new_n2821_) & (~new_n2826_ | ~new_n2821_ | ~new_n2833_ | new_n2790_ | new_n2796_ | new_n2815_ | new_n2802_ | ~new_n2809_) & (~new_n2790_ | ~new_n2821_ | ~new_n2802_ | ~new_n2809_ | new_n2826_ | ~new_n2815_ | new_n2833_);
  assign new_n2863_ = new_n2864_ & P3_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign new_n2864_ = new_n2786_ & new_n2781_ & ((P3_INSTADDRPOINTER_REG_7__SCAN_IN & (~new_n2904_ | (new_n2865_ ^ ~new_n2906_))) | (P3_INSTADDRPOINTER_REG_8__SCAN_IN & new_n2865_ & ~new_n2906_) | (~new_n2904_ & (~new_n2865_ | new_n2906_) & (new_n2865_ | ~new_n2906_))) & P3_INSTADDRPOINTER_REG_9__SCAN_IN & (P3_INSTADDRPOINTER_REG_8__SCAN_IN | (new_n2865_ & ~new_n2906_));
  assign new_n2865_ = ~new_n2899_ & ~new_n2894_ & new_n2866_ & ~new_n2889_;
  assign new_n2866_ = ~new_n2878_ & (~new_n2867_ | (~new_n2873_ & ~new_n2883_));
  assign new_n2867_ = new_n2870_ & new_n2871_ & new_n2872_ & new_n2869_ & (~new_n2804_ | ~P3_INSTQUEUE_REG_0__2__SCAN_IN) & (~new_n2868_ | ~P3_INSTQUEUE_REG_15__2__SCAN_IN);
  assign new_n2868_ = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign new_n2869_ = (~P3_INSTQUEUE_REG_5__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_9__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2870_ = (~P3_INSTQUEUE_REG_14__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_7__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_3__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2871_ = (~P3_INSTQUEUE_REG_10__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_1__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_12__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2872_ = (~P3_INSTQUEUE_REG_4__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_11__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2873_ = new_n2875_ & new_n2876_ & new_n2877_ & new_n2874_ & (~new_n2804_ | ~P3_INSTQUEUE_REG_0__1__SCAN_IN) & (~new_n2868_ | ~P3_INSTQUEUE_REG_15__1__SCAN_IN);
  assign new_n2874_ = (~P3_INSTQUEUE_REG_5__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_9__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2875_ = (~P3_INSTQUEUE_REG_14__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_7__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_3__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2876_ = (~P3_INSTQUEUE_REG_10__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_1__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_12__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2877_ = (~P3_INSTQUEUE_REG_4__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_11__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2878_ = new_n2880_ & new_n2881_ & new_n2882_ & new_n2879_ & (~new_n2803_ | ~P3_INSTQUEUE_REG_8__3__SCAN_IN) & (~new_n2868_ | ~P3_INSTQUEUE_REG_15__3__SCAN_IN);
  assign new_n2879_ = (~P3_INSTQUEUE_REG_0__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_3__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2880_ = (~P3_INSTQUEUE_REG_10__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_11__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_1__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2881_ = (~P3_INSTQUEUE_REG_14__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_5__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2882_ = (~P3_INSTQUEUE_REG_9__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_7__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2883_ = new_n2884_ & new_n2885_ & new_n2886_ & new_n2887_ & new_n2888_;
  assign new_n2884_ = (~P3_INSTQUEUE_REG_5__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_9__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2885_ = (~P3_INSTQUEUE_REG_15__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_0__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n2886_ = (~P3_INSTQUEUE_REG_14__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_7__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_3__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2887_ = (~P3_INSTQUEUE_REG_10__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_1__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_12__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2888_ = (~P3_INSTQUEUE_REG_4__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_11__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2889_ = new_n2891_ & new_n2892_ & new_n2893_ & new_n2890_ & (~new_n2803_ | ~P3_INSTQUEUE_REG_8__4__SCAN_IN) & (~new_n2868_ | ~P3_INSTQUEUE_REG_15__4__SCAN_IN);
  assign new_n2890_ = (~P3_INSTQUEUE_REG_0__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_3__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2891_ = (~P3_INSTQUEUE_REG_10__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_11__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_1__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2892_ = (~P3_INSTQUEUE_REG_14__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_5__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2893_ = (~P3_INSTQUEUE_REG_9__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_7__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2894_ = new_n2896_ & new_n2897_ & new_n2898_ & new_n2895_ & (~new_n2803_ | ~P3_INSTQUEUE_REG_8__5__SCAN_IN) & (~new_n2868_ | ~P3_INSTQUEUE_REG_15__5__SCAN_IN);
  assign new_n2895_ = (~P3_INSTQUEUE_REG_0__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_7__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_10__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2896_ = (~P3_INSTQUEUE_REG_9__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_11__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_13__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2897_ = (~P3_INSTQUEUE_REG_1__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_5__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_4__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2898_ = (~P3_INSTQUEUE_REG_14__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_3__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_6__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2899_ = new_n2901_ & new_n2902_ & new_n2903_ & new_n2900_ & (~new_n2803_ | ~P3_INSTQUEUE_REG_8__6__SCAN_IN) & (~new_n2868_ | ~P3_INSTQUEUE_REG_15__6__SCAN_IN);
  assign new_n2900_ = (~P3_INSTQUEUE_REG_0__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_7__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_10__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2901_ = (~P3_INSTQUEUE_REG_9__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_11__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_13__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2902_ = (~P3_INSTQUEUE_REG_1__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_5__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_4__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2903_ = (~P3_INSTQUEUE_REG_14__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_3__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_6__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2904_ = (~P3_INSTADDRPOINTER_REG_6__SCAN_IN | (~new_n2899_ & ~new_n2894_ & new_n2866_ & ~new_n2889_) | (new_n2899_ & (new_n2894_ | ~new_n2866_ | new_n2889_))) & ((~P3_INSTADDRPOINTER_REG_6__SCAN_IN & (new_n2899_ ^ (~new_n2894_ & new_n2866_ & ~new_n2889_))) | ((~P3_INSTADDRPOINTER_REG_5__SCAN_IN | (~new_n2894_ & new_n2866_ & ~new_n2889_) | (new_n2894_ & (~new_n2866_ | new_n2889_))) & ((~P3_INSTADDRPOINTER_REG_5__SCAN_IN & (new_n2894_ ^ (new_n2866_ & ~new_n2889_))) | (~P3_INSTADDRPOINTER_REG_4__SCAN_IN & (~new_n2866_ ^ ~new_n2889_)) | (~new_n2905_ & (~P3_INSTADDRPOINTER_REG_4__SCAN_IN | (new_n2866_ & ~new_n2889_) | (~new_n2866_ & new_n2889_))))));
  assign new_n2905_ = (P3_INSTADDRPOINTER_REG_3__SCAN_IN | (~new_n2878_ ^ (~new_n2867_ | (~new_n2873_ & ~new_n2883_)))) & ((P3_INSTADDRPOINTER_REG_3__SCAN_IN & (new_n2878_ | (new_n2867_ & (new_n2873_ | new_n2883_))) & (~new_n2878_ | ~new_n2867_ | (~new_n2873_ & ~new_n2883_))) | ((P3_INSTADDRPOINTER_REG_2__SCAN_IN | (new_n2867_ & (new_n2873_ | new_n2883_)) | (~new_n2867_ & ~new_n2873_ & ~new_n2883_)) & ((P3_INSTADDRPOINTER_REG_2__SCAN_IN & (~new_n2867_ ^ (new_n2873_ | new_n2883_))) | (((~new_n2873_ & P3_INSTADDRPOINTER_REG_1__SCAN_IN) | ~new_n2883_ | P3_INSTADDRPOINTER_REG_0__SCAN_IN) & (~new_n2873_ | P3_INSTADDRPOINTER_REG_1__SCAN_IN) & (new_n2873_ | new_n2883_)))));
  assign new_n2906_ = new_n2908_ & new_n2909_ & new_n2910_ & new_n2907_ & (~new_n2803_ | ~P3_INSTQUEUE_REG_8__7__SCAN_IN) & (~new_n2868_ | ~P3_INSTQUEUE_REG_15__7__SCAN_IN);
  assign new_n2907_ = (~P3_INSTQUEUE_REG_0__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_7__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_10__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2908_ = (~P3_INSTQUEUE_REG_9__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_11__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_13__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2909_ = (~P3_INSTQUEUE_REG_1__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_2__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_5__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_4__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n2910_ = (~P3_INSTQUEUE_REG_14__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_3__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_6__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n2911_ = new_n2912_ & P3_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign new_n2912_ = P3_INSTADDRPOINTER_REG_21__SCAN_IN & P3_INSTADDRPOINTER_REG_20__SCAN_IN & P3_INSTADDRPOINTER_REG_19__SCAN_IN & new_n2781_ & new_n2924_ & (new_n2913_ | ~new_n2922_);
  assign new_n2913_ = ~new_n2914_ & ~new_n2915_ & (~new_n2921_ | (~new_n2916_ & (new_n2918_ | ~new_n2920_) & (new_n2917_ | P3_INSTADDRPOINTER_REG_4__SCAN_IN)));
  assign new_n2914_ = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN & (new_n2906_ ^ (~new_n2899_ & ~new_n2894_ & ~new_n2889_ & ~new_n2878_ & ~new_n2867_ & ~new_n2873_));
  assign new_n2915_ = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN & (new_n2899_ ^ (~new_n2894_ & ~new_n2889_ & ~new_n2878_ & ~new_n2867_ & ~new_n2873_));
  assign new_n2916_ = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN & (new_n2894_ ^ (~new_n2889_ & ~new_n2878_ & ~new_n2867_ & ~new_n2873_));
  assign new_n2917_ = ~new_n2889_ ^ (~new_n2878_ & ~new_n2867_ & ~new_n2873_);
  assign new_n2918_ = (P3_INSTADDRPOINTER_REG_3__SCAN_IN | (~new_n2878_ ^ (~new_n2867_ & ~new_n2873_))) & (P3_INSTADDRPOINTER_REG_2__SCAN_IN | (new_n2867_ ^ new_n2873_)) & ((P3_INSTADDRPOINTER_REG_2__SCAN_IN & (~new_n2867_ | ~new_n2873_) & (new_n2867_ | new_n2873_)) | ((new_n2873_ | P3_INSTADDRPOINTER_REG_1__SCAN_IN) & (new_n2919_ | (new_n2873_ & P3_INSTADDRPOINTER_REG_1__SCAN_IN))));
  assign new_n2919_ = P3_INSTADDRPOINTER_REG_0__SCAN_IN & (~new_n2884_ | ~new_n2885_ | ~new_n2886_ | ~new_n2887_ | ~new_n2888_);
  assign new_n2920_ = (~P3_INSTADDRPOINTER_REG_4__SCAN_IN | (~new_n2889_ & ~new_n2878_ & ~new_n2867_ & ~new_n2873_) | (new_n2889_ & (new_n2878_ | new_n2867_ | new_n2873_))) & (~P3_INSTADDRPOINTER_REG_3__SCAN_IN | (~new_n2878_ & ~new_n2867_ & ~new_n2873_) | (new_n2878_ & (new_n2867_ | new_n2873_)));
  assign new_n2921_ = (~P3_INSTADDRPOINTER_REG_6__SCAN_IN | (~new_n2899_ & ~new_n2894_ & ~new_n2889_ & ~new_n2878_ & ~new_n2867_ & ~new_n2873_) | (new_n2899_ & (new_n2894_ | new_n2889_ | new_n2878_ | new_n2867_ | new_n2873_))) & (~P3_INSTADDRPOINTER_REG_5__SCAN_IN | (~new_n2894_ & ~new_n2889_ & ~new_n2878_ & ~new_n2867_ & ~new_n2873_) | (new_n2894_ & (new_n2889_ | new_n2878_ | new_n2867_ | new_n2873_)));
  assign new_n2922_ = (~P3_INSTADDRPOINTER_REG_7__SCAN_IN | (new_n2923_ & ~new_n2906_) | (~new_n2923_ & new_n2906_)) & (~P3_INSTADDRPOINTER_REG_8__SCAN_IN | ~new_n2923_ | new_n2906_);
  assign new_n2923_ = ~new_n2899_ & ~new_n2894_ & ~new_n2889_ & ~new_n2878_ & ~new_n2867_ & ~new_n2873_;
  assign new_n2924_ = P3_INSTADDRPOINTER_REG_9__SCAN_IN & (new_n2925_ | P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  assign new_n2925_ = ~new_n2906_ & ~new_n2899_ & ~new_n2894_ & ~new_n2889_ & ~new_n2878_ & ~new_n2867_ & ~new_n2873_;
  assign new_n2926_ = new_n2927_ & new_n2906_;
  assign new_n2927_ = ~new_n2802_ & ~new_n2809_ & new_n2833_ & ~new_n2790_ & ~new_n2796_ & new_n2815_ & ~new_n2826_ & ~new_n2821_;
  assign new_n2928_ = new_n2802_ & ~new_n2809_ & new_n2833_ & ~new_n2790_ & ~new_n2796_ & new_n2815_ & ~new_n2826_ & ~new_n2821_;
  assign new_n2929_ = new_n2935_ & ((((new_n2925_ & ~P3_INSTADDRPOINTER_REG_24__SCAN_IN) | (new_n2925_ & ~P3_INSTADDRPOINTER_REG_23__SCAN_IN) | ~new_n2930_ | (new_n2925_ & ~P3_INSTADDRPOINTER_REG_22__SCAN_IN)) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_24__SCAN_IN) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_23__SCAN_IN) & (new_n2925_ | new_n2936_) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_25__SCAN_IN) & (~new_n2925_ | P3_INSTADDRPOINTER_REG_25__SCAN_IN)) | ((((~new_n2925_ | P3_INSTADDRPOINTER_REG_24__SCAN_IN) & (~new_n2925_ | P3_INSTADDRPOINTER_REG_23__SCAN_IN) & new_n2930_ & (~new_n2925_ | P3_INSTADDRPOINTER_REG_22__SCAN_IN)) | (~new_n2925_ & P3_INSTADDRPOINTER_REG_24__SCAN_IN) | (~new_n2925_ & P3_INSTADDRPOINTER_REG_23__SCAN_IN) | (~new_n2925_ & ~new_n2936_) | (~new_n2925_ & P3_INSTADDRPOINTER_REG_22__SCAN_IN)) & (new_n2925_ ^ P3_INSTADDRPOINTER_REG_25__SCAN_IN)) | ((~new_n2925_ ^ ~P3_INSTADDRPOINTER_REG_23__SCAN_IN) & ((new_n2930_ & (~new_n2925_ | P3_INSTADDRPOINTER_REG_22__SCAN_IN)) | (~new_n2925_ & ~new_n2936_) | (~new_n2925_ & P3_INSTADDRPOINTER_REG_22__SCAN_IN))) | ((~new_n2925_ | P3_INSTADDRPOINTER_REG_23__SCAN_IN) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_23__SCAN_IN) & (~new_n2930_ | (new_n2925_ & ~P3_INSTADDRPOINTER_REG_22__SCAN_IN)) & (new_n2925_ | new_n2936_) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN)));
  assign new_n2930_ = (~new_n2925_ | new_n2786_) & ((~new_n2925_ & (P3_INSTADDRPOINTER_REG_17__SCAN_IN | P3_INSTADDRPOINTER_REG_16__SCAN_IN | (~new_n2925_ & P3_INSTADDRPOINTER_REG_15__SCAN_IN) | ((~new_n2925_ | P3_INSTADDRPOINTER_REG_15__SCAN_IN) & ((~new_n2925_ & P3_INSTADDRPOINTER_REG_14__SCAN_IN) | (~new_n2931_ & (~new_n2925_ | P3_INSTADDRPOINTER_REG_14__SCAN_IN)))))) | ((~new_n2925_ | P3_INSTADDRPOINTER_REG_15__SCAN_IN) & ((~new_n2925_ & P3_INSTADDRPOINTER_REG_14__SCAN_IN) | (~new_n2931_ & (~new_n2925_ | P3_INSTADDRPOINTER_REG_14__SCAN_IN))) & P3_INSTADDRPOINTER_REG_17__SCAN_IN & P3_INSTADDRPOINTER_REG_16__SCAN_IN & P3_INSTADDRPOINTER_REG_18__SCAN_IN));
  assign new_n2931_ = new_n2933_ & ((new_n2925_ & ~new_n2934_) | (new_n2925_ & ~P3_INSTADDRPOINTER_REG_11__SCAN_IN) | (new_n2925_ & ~P3_INSTADDRPOINTER_REG_10__SCAN_IN) | (~new_n2913_ & new_n2932_) | (new_n2925_ & ~new_n2784_));
  assign new_n2932_ = (~P3_INSTADDRPOINTER_REG_7__SCAN_IN | (new_n2923_ & ~new_n2906_) | (~new_n2923_ & new_n2906_)) & (~P3_INSTADDRPOINTER_REG_8__SCAN_IN | (new_n2923_ & ~new_n2906_));
  assign new_n2933_ = (new_n2925_ | ~P3_INSTADDRPOINTER_REG_11__SCAN_IN) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_9__SCAN_IN) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_10__SCAN_IN) & (new_n2925_ | (~P3_INSTADDRPOINTER_REG_12__SCAN_IN & ~P3_INSTADDRPOINTER_REG_13__SCAN_IN));
  assign new_n2934_ = P3_INSTADDRPOINTER_REG_12__SCAN_IN & P3_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign new_n2935_ = new_n2927_ & ~new_n2906_;
  assign new_n2936_ = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN & ~P3_INSTADDRPOINTER_REG_21__SCAN_IN & ~P3_INSTADDRPOINTER_REG_18__SCAN_IN & ~P3_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign new_n2937_ = new_n2950_ & ((~new_n2938_ & new_n2815_) | ~new_n2948_ | ~new_n2949_ | (new_n2942_ & new_n2947_ & ~new_n2802_ & ~new_n2815_));
  assign new_n2938_ = (new_n2802_ | ((~new_n2942_ | ~new_n2796_) & (~new_n2939_ | new_n2790_))) & (~new_n2945_ | (~new_n2809_ & (~new_n2802_ | new_n2790_ | new_n2796_))) & (~new_n2942_ | ~new_n2796_ | ~new_n2790_ | ~new_n2947_);
  assign new_n2939_ = ((~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) | (~new_n2940_ & (~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN))) & ((new_n2940_ & (~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) & (P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)) | (~new_n2940_ & (~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)) | ~new_n2941_ | (((P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & ((~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN))));
  assign new_n2940_ = (P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) & ((P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) | ((P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & ((P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) | ((P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & ((P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))))));
  assign new_n2941_ = ((~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) ^ ((P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & ((P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) | ((P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & ((P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)))))) & (((~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | ((~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))) ^ (P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN));
  assign new_n2942_ = ~new_n2943_ & ((~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) | (~new_n2940_ & (~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN))) & (~new_n2944_ | (new_n2940_ & (~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) & (P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)) | (~new_n2940_ & (~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)));
  assign new_n2943_ = READY2 & READY22_REG_SCAN_IN;
  assign new_n2944_ = ((~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) ^ ((P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & ((P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) | ((P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & ((P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)))))) & (((~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | ((~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))) ^ (P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)) & (((P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) | (P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & (~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)));
  assign new_n2945_ = ((~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) | (~new_n2940_ & (~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN))) & (~new_n2946_ | (new_n2940_ & (P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) & (~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)) | (~new_n2940_ & (P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ^ P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)));
  assign new_n2946_ = ((~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) ^ ((P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & ((P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) | ((P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & ((P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)))))) & (((P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & ((P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & (P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)) | (((~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | ((~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))) & (P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)) | ((P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)));
  assign new_n2947_ = ~P3_STATE_REG_0__SCAN_IN & (~P3_STATE_REG_2__SCAN_IN ^ ~P3_STATE_REG_1__SCAN_IN);
  assign new_n2948_ = (~new_n2802_ | new_n2809_ | ((~new_n2790_ | new_n2796_) & ~new_n2826_ & (new_n2790_ | ~new_n2796_))) & ((new_n2833_ & ~new_n2790_ & ~new_n2796_ & ~new_n2826_ & new_n2821_ & new_n2809_ & ~new_n2815_) | ((new_n2802_ | ~new_n2809_) & new_n2815_ & ~new_n2821_ & (~new_n2809_ | ~new_n2833_) & ~new_n2826_ & (new_n2790_ | ~new_n2796_) & (new_n2796_ | new_n2802_ | ~new_n2790_ | ~new_n2833_)));
  assign new_n2949_ = (~new_n2942_ | ~new_n2802_ | new_n2815_) & (~new_n2815_ | new_n2833_ | (new_n2790_ & ~new_n2796_)) & (~new_n2945_ | new_n2809_ | new_n2833_);
  assign new_n2950_ = P3_STATE2_REG_0__SCAN_IN & P3_STATE2_REG_2__SCAN_IN & ~P3_STATE2_REG_1__SCAN_IN;
  assign new_n2951_ = ((~new_n2952_ & new_n2953_) | ~new_n2505_ | ~new_n2512_ | (new_n2952_ & ~new_n2953_)) & (new_n2505_ | ~P1_EAX_REG_5__SCAN_IN) & (~new_n2505_ | new_n2512_ | (new_n2954_ ? ~BUF1_REG_5__SCAN_IN : ~DATAI_5_));
  assign new_n2952_ = (~new_n2269_ | ~new_n2271_) & ((~new_n2269_ & ~new_n2271_) | ((new_n2278_ | ~new_n2276_ | ~new_n2237_) & (~new_n2282_ | (new_n2278_ & (~new_n2276_ | ~new_n2237_)))));
  assign new_n2953_ = new_n2263_ ^ (new_n2261_ & new_n2237_);
  assign new_n2954_ = P1_ADDRESS_REG_29__SCAN_IN & (~new_n2957_ | ~new_n2958_ | ~new_n2955_ | ~new_n2956_);
  assign new_n2955_ = ~P1_ADDRESS_REG_12__SCAN_IN & ~P1_ADDRESS_REG_11__SCAN_IN & ~P1_ADDRESS_REG_14__SCAN_IN & ~P1_ADDRESS_REG_13__SCAN_IN & ~P1_ADDRESS_REG_10__SCAN_IN & ~P1_ADDRESS_REG_9__SCAN_IN & ~P1_ADDRESS_REG_8__SCAN_IN & ~P1_ADDRESS_REG_7__SCAN_IN;
  assign new_n2956_ = ~P1_ADDRESS_REG_0__SCAN_IN & ~P1_ADDRESS_REG_2__SCAN_IN & ~P1_ADDRESS_REG_1__SCAN_IN & ~P1_ADDRESS_REG_4__SCAN_IN & ~P1_ADDRESS_REG_3__SCAN_IN & ~P1_ADDRESS_REG_6__SCAN_IN & ~P1_ADDRESS_REG_5__SCAN_IN;
  assign new_n2957_ = ~P1_ADDRESS_REG_28__SCAN_IN & ~P1_ADDRESS_REG_27__SCAN_IN & ~P1_ADDRESS_REG_26__SCAN_IN & ~P1_ADDRESS_REG_25__SCAN_IN & ~P1_ADDRESS_REG_24__SCAN_IN & ~P1_ADDRESS_REG_23__SCAN_IN;
  assign new_n2958_ = ~P1_ADDRESS_REG_20__SCAN_IN & ~P1_ADDRESS_REG_19__SCAN_IN & ~P1_ADDRESS_REG_22__SCAN_IN & ~P1_ADDRESS_REG_21__SCAN_IN & ~P1_ADDRESS_REG_18__SCAN_IN & ~P1_ADDRESS_REG_17__SCAN_IN & ~P1_ADDRESS_REG_16__SCAN_IN & ~P1_ADDRESS_REG_15__SCAN_IN;
  assign new_n2959_ = new_n3051_ & new_n3072_ & new_n3079_ & new_n3096_ & new_n3028_ & new_n2999_ & ~new_n2960_ & ~new_n2983_;
  assign new_n2960_ = (new_n2961_ | ~P2_INSTQUEUE_REG_6__0__SCAN_IN) & new_n2973_ & (new_n2971_ | ~new_n2982_);
  assign new_n2961_ = new_n2965_ & ((~new_n1418_ & new_n2967_) | (~new_n2969_ & (~new_n2968_ | new_n2962_ | new_n2964_)));
  assign new_n2962_ = new_n2963_ & (~new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_));
  assign new_n2963_ = new_n1670_ & ((~new_n1315_ | ~P2_INSTQUEUE_REG_0__1__SCAN_IN) ^ (~new_n1417_ | (new_n1413_ & new_n1407_)));
  assign new_n2964_ = ~new_n1670_ & new_n1666_ & (~new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_));
  assign new_n2965_ = new_n2966_ & ((~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & new_n2967_ & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (~P2_STATE2_REG_3__SCAN_IN & (new_n1854_ | ~P2_STATE2_REG_2__SCAN_IN)));
  assign new_n2966_ = ~P2_STATE2_REG_0__SCAN_IN & ((P2_STATE2_REG_3__SCAN_IN & ~new_n1762_ & (new_n1768_ | ~new_n1781_)) | (P2_STATE2_REG_2__SCAN_IN ^ P2_STATE2_REG_1__SCAN_IN));
  assign new_n2967_ = ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n2968_ = ~P2_STATE2_REG_0__SCAN_IN & ((P2_STATE2_REG_3__SCAN_IN & ~new_n1762_ & (new_n1768_ | ~new_n1781_)) | (P2_STATE2_REG_2__SCAN_IN ^ P2_STATE2_REG_1__SCAN_IN)) & P2_STATEBS16_REG_SCAN_IN & ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN;
  assign new_n2969_ = new_n2970_ & ~P2_STATEBS16_REG_SCAN_IN;
  assign new_n2970_ = ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN;
  assign new_n2971_ = ~new_n2972_ & ((P2_STATEBS16_REG_SCAN_IN & (new_n2962_ | new_n2964_)) | ~new_n2967_ | ~new_n2970_ | new_n1418_);
  assign new_n2972_ = P2_STATE2_REG_2__SCAN_IN & (new_n1854_ | (~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & new_n2967_ & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN));
  assign new_n2973_ = (~new_n2964_ | ~new_n2968_ | ~new_n2975_) & ~new_n2974_ & (~new_n2962_ | ~new_n2968_ | ~new_n2981_);
  assign new_n2974_ = ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & new_n2967_ & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~new_n1370_ & new_n2966_ & P2_STATE2_REG_3__SCAN_IN;
  assign new_n2975_ = new_n2976_ ? BUF1_REG_16__SCAN_IN : BUF2_REG_16__SCAN_IN;
  assign new_n2976_ = P2_ADDRESS_REG_29__SCAN_IN & (~new_n2979_ | ~new_n2980_ | ~new_n2977_ | ~new_n2978_);
  assign new_n2977_ = ~P2_ADDRESS_REG_12__SCAN_IN & ~P2_ADDRESS_REG_11__SCAN_IN & ~P2_ADDRESS_REG_14__SCAN_IN & ~P2_ADDRESS_REG_13__SCAN_IN & ~P2_ADDRESS_REG_10__SCAN_IN & ~P2_ADDRESS_REG_9__SCAN_IN & ~P2_ADDRESS_REG_8__SCAN_IN & ~P2_ADDRESS_REG_7__SCAN_IN;
  assign new_n2978_ = ~P2_ADDRESS_REG_0__SCAN_IN & ~P2_ADDRESS_REG_2__SCAN_IN & ~P2_ADDRESS_REG_1__SCAN_IN & ~P2_ADDRESS_REG_4__SCAN_IN & ~P2_ADDRESS_REG_3__SCAN_IN & ~P2_ADDRESS_REG_6__SCAN_IN & ~P2_ADDRESS_REG_5__SCAN_IN;
  assign new_n2979_ = ~P2_ADDRESS_REG_28__SCAN_IN & ~P2_ADDRESS_REG_27__SCAN_IN & ~P2_ADDRESS_REG_26__SCAN_IN & ~P2_ADDRESS_REG_25__SCAN_IN & ~P2_ADDRESS_REG_24__SCAN_IN & ~P2_ADDRESS_REG_23__SCAN_IN;
  assign new_n2980_ = ~P2_ADDRESS_REG_20__SCAN_IN & ~P2_ADDRESS_REG_19__SCAN_IN & ~P2_ADDRESS_REG_22__SCAN_IN & ~P2_ADDRESS_REG_21__SCAN_IN & ~P2_ADDRESS_REG_18__SCAN_IN & ~P2_ADDRESS_REG_17__SCAN_IN & ~P2_ADDRESS_REG_16__SCAN_IN & ~P2_ADDRESS_REG_15__SCAN_IN;
  assign new_n2981_ = new_n2976_ ? BUF1_REG_24__SCAN_IN : BUF2_REG_24__SCAN_IN;
  assign new_n2982_ = new_n2966_ & (new_n2976_ ? BUF1_REG_0__SCAN_IN : BUF2_REG_0__SCAN_IN);
  assign new_n2983_ = new_n2984_ & (new_n2998_ | (new_n2996_ & ~new_n2993_ & ~new_n2995_));
  assign new_n2984_ = (P1_INSTQUEUE_REG_2__1__SCAN_IN | P1_INSTQUEUE_REG_2__6__SCAN_IN) & ~new_n2991_ & (~new_n2985_ | ~new_n2988_);
  assign new_n2985_ = ~new_n2986_ & ~new_n2987_;
  assign new_n2986_ = new_n2121_ ^ ~new_n2155_;
  assign new_n2987_ = ~new_n2122_ ^ (new_n2130_ | (P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & (new_n2127_ | ~new_n2051_ | ~new_n2128_)));
  assign new_n2988_ = ~new_n2989_ & ~new_n2990_;
  assign new_n2989_ = ~new_n2133_ ^ (~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_))));
  assign new_n2990_ = ~new_n2131_ ^ ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)));
  assign new_n2991_ = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & new_n2992_ & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n2992_ = ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n2993_ = new_n2994_ & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ ^ (new_n2148_ ^ new_n2200_));
  assign new_n2994_ = new_n2156_ ^ ~new_n2288_;
  assign new_n2995_ = ~new_n2994_ & new_n2284_ & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & (new_n2154_ ^ (new_n2148_ ^ new_n2200_));
  assign new_n2996_ = P1_STATEBS16_REG_SCAN_IN & ~P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_2__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN & (new_n2997_ | (P1_STATE2_REG_3__SCAN_IN & (new_n2478_ | new_n2482_)));
  assign new_n2997_ = P1_STATE2_REG_2__SCAN_IN ^ P1_STATE2_REG_1__SCAN_IN;
  assign new_n2998_ = new_n2576_ & ~P1_STATEBS16_REG_SCAN_IN;
  assign new_n2999_ = (~new_n3020_ | (~new_n3014_ & P1_INSTQUEUE_REG_7__2__SCAN_IN)) & (~new_n3006_ | (~new_n3000_ & P1_INSTQUEUE_REG_5__1__SCAN_IN));
  assign new_n3000_ = new_n3002_ & (new_n3005_ | (new_n3004_ & new_n2990_ & new_n2133_) | (~new_n2998_ & (new_n3001_ | ~new_n2996_)));
  assign new_n3001_ = (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ | (new_n2148_ & new_n2200_) | (~new_n2148_ & ~new_n2200_)) & (~new_n2154_ | (new_n2148_ ^ new_n2200_));
  assign new_n3002_ = new_n3003_ & ((~P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_2__SCAN_IN) | ((P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_STATE2_REG_3__SCAN_IN) & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN));
  assign new_n3003_ = ~P1_STATE2_REG_0__SCAN_IN & (new_n2997_ | (~new_n2477_ & P1_STATE2_REG_3__SCAN_IN));
  assign new_n3004_ = ~new_n2155_ & new_n2987_;
  assign new_n3005_ = P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n3006_ = (~new_n3007_ | new_n3008_) & (~new_n3011_ | ~new_n3001_ | new_n2994_) & (~new_n3013_ | ~new_n3005_) & (~new_n3012_ | ~new_n3001_ | ~new_n2994_);
  assign new_n3007_ = new_n3003_ & (new_n2954_ ? BUF1_REG_1__SCAN_IN : DATAI_1_);
  assign new_n3008_ = ~new_n3010_ & (~new_n3009_ | (P1_STATEBS16_REG_SCAN_IN & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ | (new_n2148_ & new_n2200_) | (~new_n2148_ & ~new_n2200_)) & (~new_n2154_ | (new_n2148_ ^ new_n2200_))));
  assign new_n3009_ = new_n2576_ & (new_n3005_ | (new_n2133_ & (new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_)))) & (~new_n2131_ | (~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_))) & new_n2987_ & (~new_n2050_ ^ new_n2143_)));
  assign new_n3010_ = P1_STATE2_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n3011_ = new_n2996_ & (new_n2954_ | DATAI_25_) & (~new_n2954_ | BUF1_REG_25__SCAN_IN);
  assign new_n3012_ = new_n2996_ & (new_n2954_ | DATAI_17_) & (~new_n2954_ | BUF1_REG_17__SCAN_IN);
  assign new_n3013_ = ~new_n2067_ & P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN & (new_n2997_ | (P1_STATE2_REG_3__SCAN_IN & (new_n2478_ | new_n2482_)));
  assign new_n3014_ = new_n3019_ & (~new_n3015_ | (~new_n2998_ & (new_n3018_ | ~new_n2996_)));
  assign new_n3015_ = ~new_n3017_ & (~new_n3016_ | ~new_n2990_ | ~new_n2133_);
  assign new_n3016_ = new_n2155_ & new_n2987_;
  assign new_n3017_ = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n3018_ = (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & new_n2284_ & (new_n2154_ | (new_n2148_ & new_n2200_) | (~new_n2148_ & ~new_n2200_)) & (~new_n2154_ | (new_n2148_ ^ new_n2200_));
  assign new_n3019_ = new_n3003_ & (~P1_STATE2_REG_3__SCAN_IN | (~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)) & (~P1_STATE2_REG_2__SCAN_IN | (P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN));
  assign new_n3020_ = (new_n3021_ | ~new_n3024_) & (~new_n3026_ | ~new_n3018_ | new_n2994_) & ~new_n3025_ & (~new_n3027_ | ~new_n3018_ | ~new_n2994_);
  assign new_n3021_ = ~new_n3023_ & (~new_n3022_ | (P1_STATEBS16_REG_SCAN_IN & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & new_n2284_ & (new_n2154_ | (new_n2148_ & new_n2200_) | (~new_n2148_ & ~new_n2200_)) & (~new_n2154_ | (new_n2148_ ^ new_n2200_))));
  assign new_n3022_ = new_n2576_ & (new_n3017_ | (new_n2133_ & (new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_)))) & (~new_n2131_ | (~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_))) & new_n2987_ & (~new_n2050_ | ~new_n2143_) & (new_n2050_ | new_n2143_)));
  assign new_n3023_ = P1_STATE2_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n3024_ = new_n3003_ & (new_n2954_ | DATAI_2_) & (~new_n2954_ | BUF1_REG_2__SCAN_IN);
  assign new_n3025_ = new_n3017_ & ~new_n2097_ & new_n3003_ & P1_STATE2_REG_3__SCAN_IN;
  assign new_n3026_ = new_n2996_ & (new_n2954_ | DATAI_26_) & (~new_n2954_ | BUF1_REG_26__SCAN_IN);
  assign new_n3027_ = new_n2996_ & (new_n2954_ | DATAI_18_) & (~new_n2954_ | BUF1_REG_18__SCAN_IN);
  assign new_n3028_ = (new_n3034_ | ~new_n3049_) & (new_n3029_ | ~new_n3048_) & (new_n3039_ | ~new_n3007_) & (new_n3043_ | ~P1_INSTQUEUE_REG_3__7__SCAN_IN);
  assign new_n3029_ = (~new_n3033_ | ~P1_STATE2_REG_2__SCAN_IN) & ((P1_STATEBS16_REG_SCAN_IN & (new_n3030_ | new_n3031_)) | new_n3032_ | P1_STATE2_REG_3__SCAN_IN | P1_STATE2_REG_2__SCAN_IN);
  assign new_n3030_ = new_n2994_ & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & new_n2284_ & (new_n2154_ | (new_n2148_ & new_n2200_) | (~new_n2148_ & ~new_n2200_)) & (~new_n2154_ | (new_n2148_ ^ new_n2200_));
  assign new_n3031_ = ~new_n2994_ & (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ ^ (new_n2148_ ^ new_n2200_));
  assign new_n3032_ = (~new_n2989_ | new_n2990_ | ~new_n2986_ | new_n2987_) & (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  assign new_n3033_ = (P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ^ (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)) & (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ^ P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN));
  assign new_n3034_ = ~new_n3038_ & (~new_n3036_ | (~new_n3035_ & P1_STATEBS16_REG_SCAN_IN));
  assign new_n3035_ = (~new_n2284_ | ~new_n2994_ | (~new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) | (~new_n2154_ ^ (new_n2148_ ^ new_n2200_))) & (new_n2994_ | (~new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) | new_n2284_ | (~new_n2154_ & (~new_n2148_ | ~new_n2200_) & (new_n2148_ | new_n2200_)) | (new_n2154_ & (~new_n2148_ ^ new_n2200_)));
  assign new_n3036_ = new_n2576_ & (new_n3037_ | (new_n2990_ & new_n2133_ & new_n2986_ & ~new_n2987_));
  assign new_n3037_ = P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n3038_ = P1_STATE2_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ^ P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)) & (~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  assign new_n3039_ = (~P1_STATE2_REG_2__SCAN_IN | ~new_n2120_ | ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) & ((~new_n3040_ & P1_STATEBS16_REG_SCAN_IN) | new_n3041_ | P1_STATE2_REG_3__SCAN_IN | P1_STATE2_REG_2__SCAN_IN);
  assign new_n3040_ = new_n2994_ ? ((~new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) | new_n2284_ | (~new_n2154_ & (~new_n2148_ | ~new_n2200_) & (new_n2148_ | new_n2200_)) | (new_n2154_ & (~new_n2148_ ^ new_n2200_))) : ((~new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) | ~new_n2284_ | (~new_n2154_ & (~new_n2148_ | ~new_n2200_) & (new_n2148_ | new_n2200_)) | (new_n2154_ & (~new_n2148_ ^ new_n2200_)));
  assign new_n3041_ = ~new_n3042_ & (~new_n2990_ | ~new_n2133_ | new_n2986_ | new_n2987_);
  assign new_n3042_ = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n3043_ = ~new_n3044_ & new_n3047_;
  assign new_n3044_ = new_n3045_ & (new_n2998_ | (new_n2996_ & (~new_n2284_ | (~new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) | (~new_n2154_ ^ (~new_n2148_ ^ ~new_n2200_)))));
  assign new_n3045_ = ~new_n3046_ & (~new_n2987_ | (new_n2050_ & new_n2143_) | (~new_n2050_ & ~new_n2143_) | (~new_n2133_ ^ (~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_))))) | (~new_n2131_ ^ ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))));
  assign new_n3046_ = new_n2992_ & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n3047_ = new_n3003_ & ((~P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_2__SCAN_IN) | (new_n2992_ & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_STATE2_REG_3__SCAN_IN)));
  assign new_n3048_ = new_n3003_ & (new_n2954_ | DATAI_6_) & (~new_n2954_ | BUF1_REG_6__SCAN_IN);
  assign new_n3049_ = new_n3003_ & ~new_n3050_;
  assign new_n3050_ = new_n2954_ ? ~BUF1_REG_7__SCAN_IN : ~DATAI_7_;
  assign new_n3051_ = (~new_n3052_ | (~new_n3000_ & P1_INSTQUEUE_REG_5__5__SCAN_IN)) & ((~new_n3057_ & P2_INSTQUEUE_REG_12__4__SCAN_IN) | ~new_n3068_ | (~new_n3065_ & new_n3071_));
  assign new_n3052_ = (new_n3008_ | ~new_n3053_) & (~new_n3054_ | ~new_n3001_ | new_n2994_) & (~new_n3056_ | ~new_n3005_) & (~new_n3055_ | ~new_n3001_ | ~new_n2994_);
  assign new_n3053_ = new_n3003_ & (new_n2954_ ? BUF1_REG_5__SCAN_IN : DATAI_5_);
  assign new_n3054_ = new_n2996_ & (new_n2954_ | DATAI_29_) & (~new_n2954_ | BUF1_REG_29__SCAN_IN);
  assign new_n3055_ = new_n2996_ & (new_n2954_ | DATAI_21_) & (~new_n2954_ | BUF1_REG_21__SCAN_IN);
  assign new_n3056_ = ~new_n2065_ & P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN & (new_n2997_ | (P1_STATE2_REG_3__SCAN_IN & (new_n2478_ | new_n2482_)));
  assign new_n3057_ = new_n3061_ & (new_n3064_ | (~new_n2969_ & (~new_n2968_ | new_n3058_ | new_n3060_)));
  assign new_n3058_ = new_n3059_ & (~new_n1664_ | (new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_))) & (new_n1664_ | ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ ^ (~new_n1409_ ^ new_n1421_));
  assign new_n3059_ = new_n1670_ & (~new_n1315_ | ~P2_INSTQUEUE_REG_0__1__SCAN_IN | (new_n1417_ & (~new_n1413_ | ~new_n1407_))) & ((new_n1315_ & P2_INSTQUEUE_REG_0__1__SCAN_IN) | ~new_n1417_ | (new_n1413_ & new_n1407_));
  assign new_n3060_ = ~new_n1670_ & ~new_n1666_ & (~new_n1664_ | (new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_))) & (new_n1664_ | ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_));
  assign new_n3061_ = new_n2966_ & (new_n3062_ | (~P2_STATE2_REG_3__SCAN_IN & (new_n1818_ | ~P2_STATE2_REG_2__SCAN_IN)));
  assign new_n3062_ = new_n3063_ & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n3063_ = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3064_ = P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & new_n1411_ & new_n1418_;
  assign new_n3065_ = ~new_n3066_ & (~new_n3067_ | (P2_STATEBS16_REG_SCAN_IN & (new_n3058_ | new_n3060_)));
  assign new_n3066_ = P2_STATE2_REG_2__SCAN_IN & (new_n1818_ | new_n3062_);
  assign new_n3067_ = new_n2970_ & (~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ^ (~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & (~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN));
  assign new_n3068_ = (~new_n3060_ | ~new_n3069_) & (~new_n3058_ | ~new_n3070_) & (~new_n3062_ | new_n1350_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n3069_ = new_n2968_ & (~new_n2976_ | BUF1_REG_20__SCAN_IN) & (new_n2976_ | BUF2_REG_20__SCAN_IN);
  assign new_n3070_ = new_n2968_ & (~new_n2976_ | BUF1_REG_28__SCAN_IN) & (new_n2976_ | BUF2_REG_28__SCAN_IN);
  assign new_n3071_ = new_n2966_ & (~new_n2976_ | BUF1_REG_4__SCAN_IN) & (new_n2976_ | BUF2_REG_4__SCAN_IN);
  assign new_n3072_ = ~new_n3076_ & (~new_n3077_ | ((new_n3075_ | new_n3073_ | ~new_n3074_) & new_n1758_ & (new_n3074_ | (~new_n3073_ & ~new_n3075_))));
  assign new_n3073_ = ~new_n1672_ & (~new_n1419_ ^ (~new_n1662_ & ~new_n1420_));
  assign new_n3074_ = (new_n1673_ | (new_n1662_ ^ new_n1420_)) & ((new_n1673_ & (~new_n1662_ | ~new_n1420_) & (new_n1662_ | new_n1420_)) | ((new_n1663_ | new_n1674_) & (~new_n1665_ | (new_n1663_ & new_n1674_))));
  assign new_n3075_ = new_n1672_ & (~new_n1419_ | new_n1662_ | new_n1420_) & (new_n1419_ | (~new_n1662_ & ~new_n1420_));
  assign new_n3076_ = new_n2757_ & (new_n2033_ | ~new_n1330_ | ~P2_EBX_REG_25__SCAN_IN) & ~new_n1907_ & (~new_n2033_ | (new_n1330_ & P2_EBX_REG_25__SCAN_IN));
  assign new_n3077_ = (~new_n1672_ | ~new_n1759_ | ~new_n1335_) & (new_n1759_ | ~P2_EAX_REG_5__SCAN_IN) & (new_n3078_ | new_n1784_ | ~new_n1759_ | new_n1335_);
  assign new_n3078_ = new_n2976_ ? ~BUF1_REG_5__SCAN_IN : ~BUF2_REG_5__SCAN_IN;
  assign new_n3079_ = (new_n3091_ | ~P1_INSTQUEUE_REG_11__3__SCAN_IN) & ((~new_n3080_ & P2_INSTQUEUE_REG_14__5__SCAN_IN) | ~new_n3088_ | (~new_n3087_ & new_n2966_ & ~new_n3078_));
  assign new_n3080_ = new_n3083_ & (new_n3086_ | (~new_n2969_ & (~new_n2968_ | new_n3081_ | new_n3082_)));
  assign new_n3081_ = new_n2963_ & (~new_n1664_ | (new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_))) & (new_n1664_ | ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_));
  assign new_n3082_ = ~new_n1670_ & new_n1666_ & (~new_n1664_ | (new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_))) & (new_n1664_ | ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_));
  assign new_n3083_ = new_n2966_ & (new_n3084_ | (~P2_STATE2_REG_3__SCAN_IN & (new_n1838_ | ~P2_STATE2_REG_2__SCAN_IN)));
  assign new_n3084_ = new_n3085_ & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n3085_ = P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3086_ = ~new_n1418_ & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3087_ = (~P2_STATE2_REG_2__SCAN_IN | (~new_n1838_ & ~new_n3084_)) & ((P2_STATEBS16_REG_SCAN_IN & (new_n3081_ | new_n3082_)) | ~new_n3086_ | P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_2__SCAN_IN);
  assign new_n3088_ = (~new_n2968_ | (~new_n3089_ & (~new_n3082_ | new_n3090_))) & (new_n1330_ | ~new_n3084_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n3089_ = new_n2963_ & (~new_n1664_ | (new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_))) & (new_n1664_ | ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_)) & (~new_n2976_ | BUF1_REG_29__SCAN_IN) & (new_n2976_ | BUF2_REG_29__SCAN_IN);
  assign new_n3090_ = new_n2976_ ? ~BUF1_REG_21__SCAN_IN : ~BUF2_REG_21__SCAN_IN;
  assign new_n3091_ = new_n3094_ & ((~new_n2998_ & (new_n3093_ | ~new_n2996_)) | new_n3095_ | (new_n3092_ & new_n3016_));
  assign new_n3092_ = new_n2989_ & ~new_n2990_;
  assign new_n3093_ = new_n2284_ & (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & (new_n2154_ ^ (new_n2148_ ^ new_n2200_));
  assign new_n3094_ = new_n3003_ & ((~P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_2__SCAN_IN) | ((P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_STATE2_REG_3__SCAN_IN) & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN));
  assign new_n3095_ = P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n3096_ = (new_n3091_ | ~P1_INSTQUEUE_REG_11__6__SCAN_IN) & ((~new_n3097_ & P1_INSTQUEUE_REG_9__3__SCAN_IN) | ~new_n3102_ | (~new_n3106_ & new_n3109_));
  assign new_n3097_ = ~new_n3098_ & new_n3101_;
  assign new_n3098_ = new_n3099_ & (new_n2998_ | (new_n2996_ & ((~new_n2277_ & (new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_))) | (new_n2277_ & ((~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_)))) | new_n2284_ | (~new_n2154_ ^ (~new_n2148_ ^ ~new_n2200_)))));
  assign new_n3099_ = ~new_n3100_ & (~new_n2987_ | (new_n2050_ ^ new_n2143_) | (~new_n2133_ & ~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))) | (new_n2133_ & (new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_))))) | (~new_n2131_ ^ ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))));
  assign new_n3100_ = P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n3101_ = new_n3003_ & ((~P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_2__SCAN_IN) | ((P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_STATE2_REG_3__SCAN_IN) & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN));
  assign new_n3102_ = (~new_n3031_ | ~new_n3104_) & (~new_n3103_ | ~new_n3105_) & (~new_n3100_ | new_n2091_ | ~new_n3003_ | ~P1_STATE2_REG_3__SCAN_IN);
  assign new_n3103_ = new_n2994_ & (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ ^ (new_n2148_ ^ new_n2200_));
  assign new_n3104_ = new_n2996_ & (new_n2954_ | DATAI_27_) & (~new_n2954_ | BUF1_REG_27__SCAN_IN);
  assign new_n3105_ = new_n2996_ & (new_n2954_ | DATAI_19_) & (~new_n2954_ | BUF1_REG_19__SCAN_IN);
  assign new_n3106_ = ~new_n3108_ & (~new_n3107_ | (P1_STATEBS16_REG_SCAN_IN & (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ ^ (new_n2148_ ^ new_n2200_))));
  assign new_n3107_ = new_n2576_ & (new_n3100_ | (new_n2987_ & (~new_n2050_ ^ new_n2143_) & (new_n2133_ | new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_)))) & (~new_n2133_ | (~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_))))) & (new_n2131_ ^ ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_))))));
  assign new_n3108_ = P1_STATE2_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n3109_ = new_n3003_ & (new_n2954_ ? BUF1_REG_3__SCAN_IN : DATAI_3_);
  assign new_n3110_ = new_n3111_ & new_n3116_ & new_n3157_ & new_n3196_ & new_n3202_ & new_n3180_ & ~new_n3216_ & ~new_n3220_;
  assign new_n3111_ = (new_n3087_ | ~new_n3114_) & (new_n2971_ | ~new_n3113_) & (new_n3087_ | ~new_n3115_) & (new_n3021_ | ~new_n3112_);
  assign new_n3112_ = new_n3003_ & (new_n2954_ | DATAI_4_) & (~new_n2954_ | BUF1_REG_4__SCAN_IN);
  assign new_n3113_ = new_n2966_ & (new_n2976_ ? BUF1_REG_7__SCAN_IN : BUF2_REG_7__SCAN_IN);
  assign new_n3114_ = new_n2966_ & (new_n2976_ ? BUF1_REG_2__SCAN_IN : BUF2_REG_2__SCAN_IN);
  assign new_n3115_ = new_n2966_ & (new_n2976_ ? BUF1_REG_1__SCAN_IN : BUF2_REG_1__SCAN_IN);
  assign new_n3116_ = new_n3117_ & (~new_n3103_ | new_n3153_) & (new_n3125_ | ~P2_INSTQUEUE_REG_1__3__SCAN_IN) & ~new_n3128_ & (~new_n3152_ | new_n3154_);
  assign new_n3117_ = (~new_n3031_ | new_n3118_) & (~new_n3120_ | ~new_n3124_) & (~new_n2993_ | ~new_n3055_) & (~new_n3121_ | (new_n3122_ & ~new_n3055_));
  assign new_n3118_ = ~new_n3011_ & ~new_n3119_ & (~new_n2996_ | (~new_n2954_ & ~DATAI_28_) | (new_n2954_ & ~BUF1_REG_28__SCAN_IN));
  assign new_n3119_ = new_n2996_ & (new_n2954_ | DATAI_22_) & (~new_n2954_ | BUF1_REG_22__SCAN_IN);
  assign new_n3120_ = ~new_n2994_ & (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ | (new_n2148_ & new_n2200_) | (~new_n2148_ & ~new_n2200_)) & (~new_n2154_ | (new_n2148_ ^ new_n2200_));
  assign new_n3121_ = ~new_n2994_ & (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & new_n2284_ & (new_n2154_ | (new_n2148_ & new_n2200_) | (~new_n2148_ & ~new_n2200_)) & (~new_n2154_ | (new_n2148_ ^ new_n2200_));
  assign new_n3122_ = ~new_n3011_ & (~new_n2996_ | new_n3123_);
  assign new_n3123_ = new_n2954_ ? ~BUF1_REG_16__SCAN_IN : ~DATAI_16_;
  assign new_n3124_ = new_n2996_ & (new_n2954_ ? BUF1_REG_31__SCAN_IN : DATAI_31_);
  assign new_n3125_ = (new_n3126_ | new_n3127_ | P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_2__SCAN_IN) & new_n2966_ & ((new_n3127_ & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (~P2_STATE2_REG_3__SCAN_IN & (new_n1804_ | ~P2_STATE2_REG_2__SCAN_IN)));
  assign new_n3126_ = P2_STATEBS16_REG_SCAN_IN & ~new_n1666_ & (~new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ ^ (~new_n1409_ ^ new_n1421_));
  assign new_n3127_ = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3128_ = ~new_n3129_ & new_n3149_ & (new_n3003_ | (new_n3151_ & (~new_n3147_ | (~new_n3130_ & new_n3138_))));
  assign new_n3129_ = (~new_n2284_ | (new_n2154_ & ~new_n2283_) | (~new_n2154_ & new_n2283_)) & new_n2576_ & P1_STATEBS16_REG_SCAN_IN & (new_n2284_ | (new_n2154_ ^ ~new_n2283_));
  assign new_n3130_ = (~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_FLUSH_REG_SCAN_IN | ~P1_STATE2_REG_1__SCAN_IN) & (((~new_n2989_ | new_n3137_) & ~new_n3131_ & new_n3134_) | P1_STATE2_REG_1__SCAN_IN | (new_n3131_ & ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN));
  assign new_n3131_ = (new_n2477_ | new_n3132_) & new_n3133_ & (~new_n2477_ | ~new_n2493_);
  assign new_n3132_ = ~new_n2511_ & (new_n2510_ | ((~new_n2494_ | ~new_n2509_) & (~new_n2567_ | (~new_n2509_ & ~new_n2585_))));
  assign new_n3133_ = new_n2571_ & (~new_n2097_ | new_n2067_ | ~new_n2073_) & (~new_n2508_ | new_n2510_ | ~new_n2266_ | ~new_n2067_ | ~new_n2073_);
  assign new_n3134_ = ((~new_n2493_ & ~new_n2511_) | (P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) | ((~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN))) & (~new_n2585_ | (~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ (P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN))) & (~new_n3135_ | (P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) | (~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & (~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN)));
  assign new_n3135_ = new_n3136_ & new_n2091_;
  assign new_n3136_ = new_n2067_ & new_n2073_ & new_n2097_ & ~new_n2065_ & ~new_n2053_ & ~new_n2079_ & new_n2085_;
  assign new_n3137_ = ((new_n2067_ & (new_n2091_ | (~new_n2065_ & ~new_n2053_ & ~new_n2079_ & new_n2085_)) & (~new_n2053_ | (new_n2065_ & new_n2079_)) & ((new_n2065_ & ~new_n2085_) | ~new_n2097_ | (~new_n2079_ & new_n2085_)) & (new_n2097_ | ((~new_n2065_ | new_n2085_) & new_n2079_ & (new_n2053_ | ~new_n2085_)))) | ~new_n2073_ | (new_n2079_ & ~new_n2065_ & ~new_n2067_)) & (new_n2067_ | ((new_n2091_ | (~new_n2053_ & (~new_n2065_ | new_n2085_) & (~new_n2085_ | new_n2065_ | ~new_n2079_))) & (new_n2097_ | ~new_n2085_) & (~new_n2073_ | ~new_n2097_ | ~new_n2091_))) & (~new_n2067_ | new_n2073_ | ((~new_n2065_ | new_n2085_) & ((~new_n2053_ & new_n2065_) | (~new_n2053_ & ~new_n2085_)))) & (new_n2073_ | new_n2079_ | (~new_n2065_ & new_n2085_)) & ((new_n2097_ & ~new_n2091_) | (new_n2073_ & (new_n2067_ | new_n2091_))) & (~new_n2053_ | new_n2067_) & (~new_n2073_ | ~new_n2097_ | ~new_n2091_ | new_n2085_ | ~new_n2065_ | ~new_n2053_ | ~new_n2079_) & (~new_n2067_ | ~new_n2073_ | new_n2097_ | ~new_n2091_ | new_n2065_ | ~new_n2079_ | new_n2053_ | new_n2085_) & (~new_n2091_ | new_n2097_ | ~new_n2085_ | ~new_n2065_ | ~new_n2053_ | ~new_n2079_) & (new_n2067_ | new_n2091_ | new_n2065_ | ~new_n2079_ | new_n2053_ | new_n2085_) & (~new_n2065_ | ~new_n2079_ | new_n2053_ | ~new_n2085_ | ~new_n2097_ | new_n2091_) & (~new_n2097_ | ~new_n2091_ | ~new_n2065_ | ~new_n2067_ | ~new_n2073_);
  assign new_n3138_ = ((~new_n3139_ & ~P1_STATE2_REG_1__SCAN_IN & (~new_n3131_ | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN)) | (P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P1_FLUSH_REG_SCAN_IN & P1_STATE2_REG_1__SCAN_IN) | (new_n3146_ & P1_FLUSH_REG_SCAN_IN & P1_STATE2_REG_1__SCAN_IN)) & ((~new_n3142_ & ~P1_STATE2_REG_1__SCAN_IN & (~new_n3131_ | ~new_n3145_)) | (~new_n3145_ & ~P1_FLUSH_REG_SCAN_IN & P1_STATE2_REG_1__SCAN_IN) | (~new_n3146_ & P1_FLUSH_REG_SCAN_IN & P1_STATE2_REG_1__SCAN_IN));
  assign new_n3139_ = new_n3140_ & (new_n3137_ | (~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))) | (new_n2131_ & (new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_))));
  assign new_n3140_ = new_n3141_ & ((~new_n3132_ & (new_n2478_ | new_n2482_)) | ~new_n3133_ | (new_n2493_ & ~new_n2478_ & ~new_n2482_));
  assign new_n3141_ = ((~new_n2493_ & (~new_n3136_ | new_n2091_)) | (P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ (P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN))) & (~new_n3136_ | ~new_n2091_ | (P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) | (~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & (~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN))) & (~new_n2585_ | (~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN) | (P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN));
  assign new_n3142_ = new_n3143_ & (new_n3137_ | (~new_n2987_ & (~new_n2121_ | new_n2155_) & (new_n2121_ | ~new_n2155_)));
  assign new_n3143_ = new_n3144_ & ((~new_n3132_ & (new_n2478_ | new_n2482_)) | ~new_n3133_ | (new_n2493_ & ~new_n2478_ & ~new_n2482_));
  assign new_n3144_ = (~new_n2585_ | (~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN)) & (new_n2332_ | (P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN));
  assign new_n3145_ = ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign new_n3146_ = P1_INSTADDRPOINTER_REG_0__SCAN_IN & (~P1_INSTADDRPOINTER_REG_31__SCAN_IN ^ ~P1_INSTADDRPOINTER_REG_1__SCAN_IN);
  assign new_n3147_ = (~new_n3148_ | ~new_n2599_ | new_n3131_ | P1_STATE2_REG_1__SCAN_IN) & ~P1_FLUSH_REG_SCAN_IN & (~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN | (~new_n3131_ & ~P1_STATE2_REG_1__SCAN_IN));
  assign new_n3148_ = new_n2265_ ^ (~new_n2133_ & ~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_))));
  assign new_n3149_ = ~new_n3150_ & (~new_n2998_ | (new_n2154_ & ~new_n2283_) | (~new_n2154_ & new_n2283_));
  assign new_n3150_ = (P1_STATE2_REG_3__SCAN_IN | ~P1_STATE2_REG_1__SCAN_IN) & (new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_)))) & (~new_n2131_ | (~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)));
  assign new_n3151_ = new_n2607_ & P1_STATE2_REG_0__SCAN_IN;
  assign new_n3152_ = ~new_n2994_ & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ | (new_n2148_ & new_n2200_) | (~new_n2148_ & ~new_n2200_)) & (~new_n2154_ | (new_n2148_ ^ new_n2200_));
  assign new_n3153_ = ~new_n3012_ & (~new_n2996_ | (~new_n2954_ & ~DATAI_20_) | (new_n2954_ & ~BUF1_REG_20__SCAN_IN));
  assign new_n3154_ = ~new_n3012_ & ~new_n3155_;
  assign new_n3155_ = new_n2996_ & ~new_n3156_;
  assign new_n3156_ = new_n2954_ ? ~BUF1_REG_23__SCAN_IN : ~DATAI_23_;
  assign new_n3157_ = new_n3160_ & new_n3163_ & (new_n3158_ | ~new_n3115_) & (~new_n3161_ | ~new_n3054_) & (new_n3167_ | new_n3176_);
  assign new_n3158_ = (~P2_STATE2_REG_2__SCAN_IN | (~new_n1806_ & (~new_n3063_ | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))) & ((new_n3159_ & P2_STATEBS16_REG_SCAN_IN) | ~new_n3063_ | P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_2__SCAN_IN);
  assign new_n3159_ = ~new_n1666_ & (~new_n1664_ | (new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_))) & (new_n1664_ | ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_));
  assign new_n3160_ = (new_n3154_ | ~new_n3161_) & (~new_n3162_ | ((new_n1665_ | (~new_n1663_ & ~new_n1674_) | (new_n1663_ & new_n1674_)) & new_n1758_ & (~new_n1665_ | (~new_n1663_ ^ ~new_n1674_))));
  assign new_n3161_ = ~new_n2994_ & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ ^ (new_n2148_ ^ new_n2200_));
  assign new_n3162_ = ((new_n2976_ ? ~BUF1_REG_3__SCAN_IN : ~BUF2_REG_3__SCAN_IN) | new_n1784_ | ~new_n1759_ | new_n1335_) & (new_n1759_ | ~P2_EAX_REG_3__SCAN_IN) & (~new_n1674_ | ~new_n1759_ | ~new_n1335_);
  assign new_n3163_ = ~new_n3164_ & (~new_n3166_ | ((~P2_STATE2_REG_2__SCAN_IN | (~new_n1804_ & (~new_n3127_ | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))) & (new_n3126_ | ~new_n3127_ | P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_2__SCAN_IN)));
  assign new_n3164_ = (new_n3011_ | new_n3165_) & new_n2994_ & (new_n2277_ ^ ((new_n2154_ | (new_n2148_ & new_n2200_)) & (new_n2148_ | new_n2200_))) & ~new_n2284_ & (new_n2154_ ^ (new_n2148_ ^ new_n2200_));
  assign new_n3165_ = new_n2996_ & (new_n2954_ | DATAI_30_) & (~new_n2954_ | BUF1_REG_30__SCAN_IN);
  assign new_n3166_ = new_n2966_ & (new_n2976_ ? BUF1_REG_3__SCAN_IN : BUF2_REG_3__SCAN_IN);
  assign new_n3167_ = ~new_n3168_ & (new_n3170_ | P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_1__SCAN_IN) & (~new_n1670_ | ~new_n3169_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n3168_ = (~new_n2727_ | ~P2_INSTADDRPOINTER_REG_0__SCAN_IN) & P2_STATE2_REG_1__SCAN_IN & (new_n2727_ | (~P2_STATE2_REG_0__SCAN_IN & ~P2_PHYADDRPOINTER_REG_0__SCAN_IN) | (P2_STATE2_REG_0__SCAN_IN & ~P2_INSTADDRPOINTER_REG_0__SCAN_IN));
  assign new_n3169_ = ~new_n1762_ & (new_n1768_ | ~new_n1781_);
  assign new_n3170_ = new_n3173_ & (new_n3171_ | (~new_n1390_ & (~new_n1328_ | ~new_n1388_) & (new_n1391_ | ~new_n1392_)) | ((new_n1390_ | (new_n1328_ & new_n1388_)) & ~new_n1391_ & new_n1392_));
  assign new_n3171_ = ~new_n2708_ & new_n3172_;
  assign new_n3172_ = (new_n1345_ | ((new_n1322_ | (((~new_n1330_ ^ new_n1317_) | (~new_n1330_ & ~new_n1350_)) & ~new_n1335_ & (new_n1350_ | (~new_n1330_ & new_n1317_)))) & new_n1367_ & (~new_n1322_ | new_n1370_ | (~new_n1335_ & (new_n1330_ | ~new_n1317_) & (~new_n1330_ | new_n1317_))))) & (~new_n1322_ | ~new_n1370_ | ((new_n1367_ | (~new_n1335_ & ~new_n1317_ & ~new_n1330_ & new_n1350_)) & (new_n1350_ ? (~new_n1317_ | ~new_n1367_) : ~new_n1335_) & ((~new_n1330_ & new_n1317_) | (new_n1345_ & (new_n1330_ | ~new_n1367_))))) & (~new_n1345_ | ~new_n1367_ | ((new_n1322_ | ~new_n1370_) & (~new_n1322_ | new_n1370_) & ((new_n1330_ & ~new_n1317_ & new_n1335_ & new_n1350_) | (new_n1322_ & (new_n1330_ | ~new_n1317_))))) & (~new_n1322_ | ~new_n1370_ | ~new_n1345_ | ~new_n1367_ | ~new_n1330_ | new_n1317_ | ~new_n1335_ | ~new_n1350_) & (new_n1350_ | (new_n1322_ & new_n1370_) | (~new_n1322_ & ~new_n1370_)) & (new_n1322_ | ~new_n1370_ | (~new_n1330_ & ~new_n1335_)) & (new_n1367_ | (~new_n1317_ & new_n1370_));
  assign new_n3173_ = (new_n3174_ | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (new_n3175_ | ~new_n1367_ | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3174_ = (new_n1335_ | new_n1317_ | new_n1330_ | ~new_n1350_ | ~new_n1370_ | ~new_n1345_ | new_n1367_) & (~new_n1345_ | ~new_n1367_ | ~new_n1330_ | new_n1335_ | ~new_n1322_ | new_n1317_ | ~new_n1370_) & (new_n1370_ | ~new_n1350_ | new_n1335_ | new_n1345_ | ~new_n1330_ | ~new_n1317_ | ~new_n1367_);
  assign new_n3175_ = ((new_n1322_ ^ new_n1370_) | new_n1335_ | new_n1350_ | new_n1345_ | new_n1330_ | ~new_n1317_) & (~new_n1330_ | ~new_n1345_ | ((~new_n1330_ | new_n1317_ | ~new_n1335_ | ~new_n1350_ | new_n1322_ | new_n1370_) & (new_n1335_ | new_n1350_ | ~new_n1317_ | ~new_n1322_ | ~new_n1370_)));
  assign new_n3176_ = ((~new_n3177_ & new_n3178_) | ~P2_STATE2_REG_0__SCAN_IN | ~P2_STATE2_REG_2__SCAN_IN | P2_STATE2_REG_1__SCAN_IN) & (P2_STATE2_REG_0__SCAN_IN ? (~P2_FLUSH_REG_SCAN_IN | ~P2_STATE2_REG_2__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN) : ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n3177_ = new_n2670_ & ~new_n1790_ & new_n2667_ & ~new_n1762_ & (new_n1768_ | ~new_n1781_);
  assign new_n3178_ = ~new_n1785_ & (~new_n1783_ | new_n1762_ | (~new_n1768_ & new_n1781_)) & new_n3179_ & (~new_n2684_ | (~new_n1762_ & (new_n1768_ | ~new_n1781_)));
  assign new_n3179_ = new_n2711_ & (~new_n1787_ | ~new_n1788_ | ~new_n2670_ | new_n1790_);
  assign new_n3180_ = (new_n3185_ | ~new_n3186_ | (~new_n3181_ & P2_INSTQUEUE_REG_15__2__SCAN_IN)) & (new_n3190_ | ~new_n3192_ | (~new_n3181_ & P2_INSTQUEUE_REG_15__6__SCAN_IN));
  assign new_n3181_ = new_n3183_ & (new_n3085_ | (~new_n2969_ & (new_n3182_ | ~new_n2968_)));
  assign new_n3182_ = new_n1666_ & (~new_n1664_ | (new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_))) & (new_n1664_ | ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_));
  assign new_n3183_ = new_n2966_ & (new_n3184_ | (~P2_STATE2_REG_3__SCAN_IN & (new_n1817_ | ~P2_STATE2_REG_2__SCAN_IN)));
  assign new_n3184_ = P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3185_ = new_n3114_ & ((P2_STATE2_REG_2__SCAN_IN & (new_n1817_ | new_n3184_)) | ((~new_n3182_ | ~P2_STATEBS16_REG_SCAN_IN) & new_n3085_ & ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN));
  assign new_n3186_ = (~new_n3082_ | ~new_n3188_) & (~new_n3187_ | ~new_n3189_) & (~new_n3184_ | new_n1367_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n3187_ = new_n3059_ & (~new_n1664_ | (new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_))) & (new_n1664_ | ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_));
  assign new_n3188_ = new_n2968_ & (new_n2976_ ? BUF1_REG_26__SCAN_IN : BUF2_REG_26__SCAN_IN);
  assign new_n3189_ = new_n2968_ & (~new_n2976_ | BUF1_REG_18__SCAN_IN) & (new_n2976_ | BUF2_REG_18__SCAN_IN);
  assign new_n3190_ = new_n3191_ & ((P2_STATE2_REG_2__SCAN_IN & (new_n1817_ | new_n3184_)) | ((~new_n3182_ | ~P2_STATEBS16_REG_SCAN_IN) & new_n3085_ & ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN));
  assign new_n3191_ = new_n2966_ & (new_n2976_ ? BUF1_REG_6__SCAN_IN : BUF2_REG_6__SCAN_IN);
  assign new_n3192_ = (~new_n3082_ | ~new_n3193_) & (~new_n3187_ | ~new_n3195_) & (~new_n3184_ | new_n1317_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n3193_ = new_n2968_ & ~new_n3194_;
  assign new_n3194_ = new_n2976_ ? ~BUF1_REG_30__SCAN_IN : ~BUF2_REG_30__SCAN_IN;
  assign new_n3195_ = new_n2968_ & (new_n2976_ ? BUF1_REG_22__SCAN_IN : BUF2_REG_22__SCAN_IN);
  assign new_n3196_ = (new_n3197_ | ~new_n3198_ | (~new_n3125_ & P2_INSTQUEUE_REG_1__4__SCAN_IN)) & (new_n3106_ | (~new_n3007_ & ~new_n3112_));
  assign new_n3197_ = new_n3071_ & ((P2_STATE2_REG_2__SCAN_IN & (new_n1804_ | (new_n3127_ & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))) | (~new_n3126_ & new_n3127_ & ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN));
  assign new_n3198_ = (~new_n3199_ | ~new_n3070_) & ~new_n3200_ & (~new_n3201_ | new_n1350_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n3199_ = ~new_n1670_ & ~new_n1666_ & (~new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ ^ (~new_n1409_ ^ new_n1421_));
  assign new_n3200_ = new_n3069_ & new_n2963_ & (~new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ ^ (~new_n1409_ ^ new_n1421_));
  assign new_n3201_ = new_n3127_ & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n3202_ = (~new_n3049_ | new_n3212_) & (new_n3203_ | ~new_n3208_ | (~new_n3207_ & new_n3166_));
  assign new_n3203_ = P2_INSTQUEUE_REG_7__3__SCAN_IN & (~new_n3205_ | (~new_n3204_ & new_n2970_ & (~new_n2967_ | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)));
  assign new_n3204_ = P2_STATEBS16_REG_SCAN_IN & new_n1666_ & (~new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_));
  assign new_n3205_ = new_n2966_ & (new_n3206_ | (~P2_STATE2_REG_3__SCAN_IN & (new_n1805_ | ~P2_STATE2_REG_2__SCAN_IN)));
  assign new_n3206_ = ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n3207_ = (~P2_STATE2_REG_2__SCAN_IN | (~new_n1805_ & ~new_n3206_)) & (new_n3204_ | ~new_n2967_ | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_2__SCAN_IN);
  assign new_n3208_ = (~new_n2964_ | ~new_n3211_) & ~new_n3209_ & (~new_n3206_ | new_n1345_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n3209_ = new_n2968_ & new_n3210_ & new_n3059_ & (~new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_));
  assign new_n3210_ = new_n2976_ ? BUF1_REG_19__SCAN_IN : BUF2_REG_19__SCAN_IN;
  assign new_n3211_ = new_n2968_ & (~new_n2976_ | BUF1_REG_27__SCAN_IN) & (new_n2976_ | BUF2_REG_27__SCAN_IN);
  assign new_n3212_ = ~new_n3215_ & (~new_n3213_ | (P1_STATEBS16_REG_SCAN_IN & (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ | (new_n2148_ & new_n2200_) | (~new_n2148_ & ~new_n2200_)) & (~new_n2154_ | (new_n2148_ ^ new_n2200_))));
  assign new_n3213_ = new_n2576_ & (new_n3214_ | (new_n2987_ & (~new_n2050_ ^ new_n2143_) & ~new_n2133_ & (new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_)))) & (~new_n2131_ | (~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))));
  assign new_n3214_ = P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n3215_ = P1_STATE2_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n3216_ = new_n3053_ & (new_n3218_ | ((~new_n3217_ | ~P1_STATEBS16_REG_SCAN_IN) & new_n2576_ & (new_n3219_ | (new_n2988_ & new_n3004_))));
  assign new_n3217_ = (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ ^ (new_n2148_ ^ new_n2200_));
  assign new_n3218_ = ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & new_n2992_ & P1_STATE2_REG_2__SCAN_IN;
  assign new_n3219_ = new_n2992_ & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n3220_ = new_n3007_ & ~new_n3221_;
  assign new_n3221_ = ~new_n3224_ & (~new_n3222_ | (P1_STATEBS16_REG_SCAN_IN & (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & new_n2284_ & (new_n2154_ | (new_n2148_ & new_n2200_) | (~new_n2148_ & ~new_n2200_)) & (~new_n2154_ | (new_n2148_ ^ new_n2200_))));
  assign new_n3222_ = new_n2576_ & (new_n3223_ | (new_n2987_ & (~new_n2050_ | ~new_n2143_) & (new_n2050_ | new_n2143_) & ~new_n2133_ & (new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_)))) & (~new_n2131_ | (~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))));
  assign new_n3223_ = P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n3224_ = P1_STATE2_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n3225_ = new_n3226_ & new_n3263_ & new_n3367_ & new_n3387_ & new_n3399_ & new_n4089_ & new_n4100_ & new_n4118_;
  assign new_n3226_ = new_n3256_ & new_n3227_ & new_n3249_ & ~new_n3261_ & (new_n3246_ | ~P2_INSTQUEUE_REG_13__1__SCAN_IN);
  assign new_n3227_ = new_n3228_ & ~new_n3232_ & ((P2_INSTQUEUE_REG_5__1__SCAN_IN & (new_n3233_ | ~new_n3235_)) | new_n3237_ | new_n3240_ | ~new_n3243_);
  assign new_n3228_ = (~new_n3229_ | new_n2994_ | ~new_n2284_ | (~new_n2277_ ^ ((new_n2154_ | (new_n2148_ & new_n2200_)) & (new_n2148_ | new_n2200_))) | (~new_n2154_ ^ (new_n2148_ ^ new_n2200_))) & (new_n3231_ | new_n2994_ | ~new_n2284_ | (~new_n2277_ ^ ((new_n2154_ | (new_n2148_ & new_n2200_)) & (new_n2148_ | new_n2200_))) | (~new_n2154_ ^ (new_n2148_ ^ new_n2200_)));
  assign new_n3229_ = new_n2996_ & ~new_n3230_;
  assign new_n3230_ = new_n2954_ ? ~BUF1_REG_24__SCAN_IN : ~DATAI_24_;
  assign new_n3231_ = (~new_n2996_ | (new_n2954_ & ~BUF1_REG_17__SCAN_IN) | (~new_n2954_ & ~DATAI_17_)) & (~new_n2996_ | (new_n2954_ & ~BUF1_REG_22__SCAN_IN) | (~new_n2954_ & ~DATAI_22_));
  assign new_n3232_ = (new_n3104_ | new_n3124_) & ~new_n2994_ & new_n2284_ & (new_n2277_ ^ ((new_n2154_ | (new_n2148_ & new_n2200_)) & (new_n2148_ | new_n2200_))) & (new_n2154_ ^ (new_n2148_ ^ new_n2200_));
  assign new_n3233_ = (~new_n3234_ | (new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) | (~new_n1412_ & (new_n1409_ | ~new_n1421_) & (~new_n1409_ | new_n1421_)) | (new_n1412_ & (new_n1409_ ^ new_n1421_))) & new_n2970_ & (~new_n2967_ | P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  assign new_n3234_ = P2_STATEBS16_REG_SCAN_IN & (new_n1414_ ^ ((~new_n1315_ | ~P2_INSTQUEUE_REG_0__1__SCAN_IN) ^ (~new_n1417_ | (new_n1413_ & new_n1407_))));
  assign new_n3235_ = new_n2966_ & (new_n3236_ | (~P2_STATE2_REG_3__SCAN_IN & (new_n1811_ | ~P2_STATE2_REG_2__SCAN_IN)));
  assign new_n3236_ = P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & new_n2967_ & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n3237_ = new_n3115_ & (new_n3238_ | (new_n3239_ & (~new_n3234_ | (new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) | (~new_n1412_ & (~new_n1409_ | new_n1421_) & (new_n1409_ | ~new_n1421_)) | (new_n1412_ & (~new_n1409_ ^ ~new_n1421_)))));
  assign new_n3238_ = P2_STATE2_REG_2__SCAN_IN & (new_n3236_ | (~new_n1413_ & new_n1803_ & (~new_n1327_ ^ (new_n1383_ | (~new_n1386_ & ~new_n1387_))) & (new_n1387_ | new_n1383_ | new_n1386_) & (~new_n1387_ | (~new_n1383_ & ~new_n1386_))));
  assign new_n3239_ = new_n2970_ & new_n2967_ & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n3240_ = new_n3241_ & new_n3242_ & (~new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_));
  assign new_n3241_ = new_n2968_ & (~new_n2976_ | BUF1_REG_25__SCAN_IN) & (new_n2976_ | BUF2_REG_25__SCAN_IN);
  assign new_n3242_ = ~new_n1670_ & (new_n1414_ ^ ((~new_n1315_ | ~P2_INSTQUEUE_REG_0__1__SCAN_IN) ^ (~new_n1417_ | (new_n1413_ & new_n1407_))));
  assign new_n3243_ = ~new_n3245_ & (~new_n3244_ | ~new_n2963_ | (new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) | (~new_n1412_ & (~new_n1409_ | new_n1421_) & (new_n1409_ | ~new_n1421_)) | (new_n1412_ & (~new_n1409_ ^ ~new_n1421_)));
  assign new_n3244_ = new_n2968_ & (new_n2976_ ? BUF1_REG_17__SCAN_IN : BUF2_REG_17__SCAN_IN);
  assign new_n3245_ = new_n3236_ & ~new_n1322_ & new_n2966_ & P2_STATE2_REG_3__SCAN_IN;
  assign new_n3246_ = new_n3247_ & (new_n3063_ | (~new_n2969_ & (new_n3159_ | ~new_n2968_)));
  assign new_n3247_ = new_n2966_ & (new_n3248_ | (~P2_STATE2_REG_3__SCAN_IN & (new_n1806_ | ~P2_STATE2_REG_2__SCAN_IN)));
  assign new_n3248_ = new_n3063_ & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n3249_ = (new_n3250_ | new_n3176_) & ((~new_n1977_ & new_n1993_) | ~new_n2691_ | (new_n1977_ & ~new_n1993_));
  assign new_n3250_ = (new_n3251_ | ~P2_STATE2_REG_1__SCAN_IN) & (~new_n3169_ | ~P2_STATE2_REG_3__SCAN_IN | (~new_n1412_ & (new_n1409_ | ~new_n1421_) & (~new_n1409_ | new_n1421_)) | (new_n1412_ & (new_n1409_ ^ new_n1421_))) & (new_n3252_ | P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_1__SCAN_IN);
  assign new_n3251_ = (~P2_INSTADDRPOINTER_REG_1__SCAN_IN | ~new_n2727_ | ~P2_INSTADDRPOINTER_REG_0__SCAN_IN) & ((P2_STATE2_REG_0__SCAN_IN ? P2_INSTADDRPOINTER_REG_1__SCAN_IN : ~P2_PHYADDRPOINTER_REG_1__SCAN_IN) | new_n2727_ | (P2_STATE2_REG_0__SCAN_IN & ~P2_INSTADDRPOINTER_REG_0__SCAN_IN) | (~P2_STATE2_REG_0__SCAN_IN & ~P2_PHYADDRPOINTER_REG_0__SCAN_IN));
  assign new_n3252_ = new_n3253_ & (new_n3171_ | (new_n1387_ & ~new_n1410_) | (~new_n1387_ & new_n1410_));
  assign new_n3253_ = (new_n3174_ | (P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN)) & (~new_n3254_ | (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) | (P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN))) & (new_n3255_ | ((~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN))));
  assign new_n3254_ = new_n1367_ & ~new_n1335_ & ~new_n1350_ & new_n1784_ & ~new_n1345_ & (~new_n1322_ ^ new_n1370_);
  assign new_n3255_ = ~new_n1375_ & (~new_n1764_ | ~new_n1761_ | ~new_n1359_);
  assign new_n3256_ = ~new_n3260_ & (~P1_INSTQUEUE_REG_15__1__SCAN_IN | (new_n3259_ & (~new_n3258_ | (~new_n2998_ & (~new_n2996_ | (new_n2276_ & new_n3257_))))));
  assign new_n3257_ = new_n2284_ & (~new_n2154_ | new_n2283_) & (new_n2154_ | ~new_n2283_);
  assign new_n3258_ = ~new_n3223_ & (~new_n3016_ | ~new_n2990_ | new_n2133_);
  assign new_n3259_ = new_n3003_ & (~P1_STATE2_REG_3__SCAN_IN | (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)) & (~P1_STATE2_REG_2__SCAN_IN | (P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN));
  assign new_n3260_ = new_n2678_ & (new_n1619_ | ~new_n1531_ | new_n1618_) & (~new_n1619_ | (new_n1531_ & ~new_n1618_));
  assign new_n3261_ = (~new_n2476_ | new_n2053_ | (new_n2287_ ^ (new_n2285_ ^ (~new_n2284_ | ~new_n2237_)))) & (new_n2476_ | ~P1_EBX_REG_1__SCAN_IN) & (~new_n3262_ | ~new_n2476_ | ~new_n2053_);
  assign new_n3262_ = ((~P1_EBX_REG_0__SCAN_IN & (~P1_INSTADDRPOINTER_REG_0__SCAN_IN | (~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_))) ? (~new_n2067_ & ~new_n2091_) : (~new_n2073_ & new_n2091_)) ^ (((new_n2067_ | new_n2073_) & (new_n2073_ | ~new_n2116_)) ^ ((new_n2067_ | new_n2091_) ^ ((~P1_EBX_REG_1__SCAN_IN | (new_n2091_ ? new_n2073_ : new_n2067_)) & (~P1_INSTADDRPOINTER_REG_1__SCAN_IN | (~new_n2067_ & ~new_n2073_) | (~new_n2073_ & new_n2116_)))));
  assign new_n3263_ = new_n3264_ & new_n3272_ & new_n3275_ & new_n3361_ & new_n3365_ & (new_n3362_ | ~P2_INSTQUEUE_REG_11__3__SCAN_IN);
  assign new_n3264_ = new_n3267_ & (~new_n3265_ | ~new_n3011_) & (~new_n3266_ | ~new_n2996_ | (~new_n2954_ & ~DATAI_28_) | (new_n2954_ & ~BUF1_REG_28__SCAN_IN));
  assign new_n3265_ = new_n2994_ & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ | (new_n2148_ & new_n2200_) | (~new_n2148_ & ~new_n2200_)) & (~new_n2154_ | (new_n2148_ ^ new_n2200_));
  assign new_n3266_ = ~new_n2994_ & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & new_n2284_ & (new_n2154_ | (new_n2148_ & new_n2200_) | (~new_n2148_ & ~new_n2200_)) & (~new_n2154_ | (new_n2148_ ^ new_n2200_));
  assign new_n3267_ = (new_n3269_ | ~new_n3268_ | (~new_n2277_ & (new_n2154_ | (new_n2148_ & new_n2200_)) & (new_n2148_ | new_n2200_)) | (new_n2277_ & ((~new_n2154_ & (~new_n2148_ | ~new_n2200_)) | (~new_n2148_ & ~new_n2200_))) | (~new_n2154_ ^ (new_n2148_ ^ new_n2200_))) & ((new_n3270_ & new_n3271_) | ~new_n3268_ | (~new_n2277_ ^ ((new_n2154_ | (new_n2148_ & new_n2200_)) & (new_n2148_ | new_n2200_))) | (~new_n2154_ ^ (new_n2148_ ^ new_n2200_)));
  assign new_n3268_ = (new_n2163_ | (~new_n2156_ & ~new_n2176_) | (~new_n2175_ ^ (new_n2169_ | (~P1_STATE2_REG_0__SCAN_IN & (~new_n2121_ ^ ~new_n2155_))))) & ((~new_n2175_ & (new_n2169_ | (~P1_STATE2_REG_0__SCAN_IN & (~new_n2121_ ^ ~new_n2155_)))) | (~new_n2163_ & (new_n2156_ | new_n2176_)) | (new_n2175_ & ~new_n2169_ & (P1_STATE2_REG_0__SCAN_IN | (new_n2121_ ^ ~new_n2155_)))) & (~new_n2156_ | (~new_n2163_ & ~new_n2176_)) & (new_n2156_ | new_n2163_ | new_n2176_);
  assign new_n3269_ = (~new_n2996_ | (new_n2954_ & ~BUF1_REG_19__SCAN_IN) | (~new_n2954_ & ~DATAI_19_)) & (~new_n2996_ | (new_n2954_ & ~BUF1_REG_22__SCAN_IN) | (~new_n2954_ & ~DATAI_22_));
  assign new_n3270_ = (~new_n2996_ | (new_n2954_ & ~BUF1_REG_25__SCAN_IN) | (~new_n2954_ & ~DATAI_25_)) & (~new_n2996_ | (new_n2954_ ? ~BUF1_REG_31__SCAN_IN : ~DATAI_31_));
  assign new_n3271_ = (~new_n2996_ | (~new_n2954_ & ~DATAI_19_) | (new_n2954_ & ~BUF1_REG_19__SCAN_IN)) & (~new_n2996_ | new_n3123_) & (~new_n2996_ | new_n3156_);
  assign new_n3272_ = (~new_n3273_ | ~new_n3211_) & (~new_n3060_ | ~new_n2968_ | ~new_n2975_) & (~new_n3273_ | ~new_n3195_) & (~new_n2964_ | ~new_n2968_ | ~new_n3274_);
  assign new_n3273_ = ~new_n1670_ & new_n1666_ & (~new_n1664_ | (new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_))) & (new_n1664_ | ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ ^ (~new_n1409_ ^ new_n1421_));
  assign new_n3274_ = new_n2976_ ? BUF1_REG_23__SCAN_IN : BUF2_REG_23__SCAN_IN;
  assign new_n3275_ = new_n3276_ & new_n3355_ & new_n3320_ & new_n3310_ & new_n3316_ & new_n3340_ & new_n3325_ & new_n3335_;
  assign new_n3276_ = ~new_n3277_ & (new_n3309_ | (~new_n2641_ & ~new_n2642_)) & ~new_n3308_ & (new_n3288_ | ~new_n3290_);
  assign new_n3277_ = new_n3281_ & (~new_n2937_ | (((~new_n3278_ & ~P3_INSTADDRPOINTER_REG_10__SCAN_IN) | ~new_n2928_ | (new_n3278_ & P3_INSTADDRPOINTER_REG_10__SCAN_IN)) & ~new_n3279_ & ~new_n3280_ & new_n3285_));
  assign new_n3278_ = ((P3_INSTADDRPOINTER_REG_7__SCAN_IN & (~new_n2904_ | (new_n2865_ ^ ~new_n2906_))) | (P3_INSTADDRPOINTER_REG_8__SCAN_IN & new_n2865_ & ~new_n2906_) | (~new_n2904_ & (~new_n2865_ | new_n2906_) & (new_n2865_ | ~new_n2906_))) & P3_INSTADDRPOINTER_REG_9__SCAN_IN & (P3_INSTADDRPOINTER_REG_8__SCAN_IN | (new_n2865_ & ~new_n2906_));
  assign new_n3279_ = ((new_n2925_ ^ ~P3_INSTADDRPOINTER_REG_10__SCAN_IN) | (~new_n2925_ & P3_INSTADDRPOINTER_REG_9__SCAN_IN) | ((new_n2913_ | ~new_n2932_) & (~new_n2925_ | (P3_INSTADDRPOINTER_REG_8__SCAN_IN & P3_INSTADDRPOINTER_REG_9__SCAN_IN)))) & new_n2935_ & ((new_n2925_ & ~P3_INSTADDRPOINTER_REG_10__SCAN_IN) | (~new_n2925_ & P3_INSTADDRPOINTER_REG_10__SCAN_IN) | ((new_n2925_ | ~P3_INSTADDRPOINTER_REG_9__SCAN_IN) & ((~new_n2913_ & new_n2932_) | (new_n2925_ & (~P3_INSTADDRPOINTER_REG_8__SCAN_IN | ~P3_INSTADDRPOINTER_REG_9__SCAN_IN)))));
  assign new_n3280_ = (P3_INSTADDRPOINTER_REG_10__SCAN_IN | (new_n2924_ & (new_n2913_ | ~new_n2922_))) & new_n2926_ & (~P3_INSTADDRPOINTER_REG_10__SCAN_IN | ~new_n2924_ | (~new_n2913_ & new_n2922_));
  assign new_n3281_ = (~P3_INSTADDRPOINTER_REG_10__SCAN_IN | new_n2937_ | new_n3282_) & (~P3_REIP_REG_10__SCAN_IN | P3_STATE2_REG_2__SCAN_IN | (~new_n2937_ & ~new_n3282_));
  assign new_n3282_ = new_n3283_ & new_n3284_;
  assign new_n3283_ = ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN;
  assign new_n3284_ = ~P3_STATE2_REG_2__SCAN_IN & ~P3_STATE2_REG_1__SCAN_IN;
  assign new_n3285_ = (new_n3286_ | (~P3_INSTADDRPOINTER_REG_10__SCAN_IN & (~new_n2783_ | ~P3_INSTADDRPOINTER_REG_2__SCAN_IN | ~P3_INSTADDRPOINTER_REG_0__SCAN_IN | ~P3_INSTADDRPOINTER_REG_1__SCAN_IN)) | (P3_INSTADDRPOINTER_REG_10__SCAN_IN & new_n2783_ & P3_INSTADDRPOINTER_REG_2__SCAN_IN & P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN)) & (~new_n2850_ | (~P3_INSTADDRPOINTER_REG_10__SCAN_IN & (~new_n2783_ | (~P3_INSTADDRPOINTER_REG_2__SCAN_IN & (~P3_INSTADDRPOINTER_REG_0__SCAN_IN | ~P3_INSTADDRPOINTER_REG_1__SCAN_IN)))) | (P3_INSTADDRPOINTER_REG_10__SCAN_IN & new_n2783_ & (P3_INSTADDRPOINTER_REG_2__SCAN_IN | (P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN)))) & (new_n3287_ | (~P3_INSTADDRPOINTER_REG_10__SCAN_IN & (~new_n2783_ | ~P3_INSTADDRPOINTER_REG_1__SCAN_IN | ~P3_INSTADDRPOINTER_REG_2__SCAN_IN)) | (P3_INSTADDRPOINTER_REG_10__SCAN_IN & new_n2783_ & P3_INSTADDRPOINTER_REG_1__SCAN_IN & P3_INSTADDRPOINTER_REG_2__SCAN_IN));
  assign new_n3286_ = (~new_n2815_ | ((~new_n2802_ | new_n2809_ | (~new_n2821_ & (~new_n2790_ | new_n2796_) & ~new_n2826_ & (new_n2790_ | ~new_n2796_))) & (~new_n2809_ | ((~new_n2790_ | ~new_n2833_) & (~new_n2802_ | new_n2790_ | new_n2796_))) & ((new_n2796_ & new_n2826_) | new_n2802_ | (~new_n2826_ & ~new_n2821_)))) & (new_n2796_ | ~new_n2821_ | (new_n2809_ & (~new_n2802_ | ~new_n2826_))) & (new_n2796_ | new_n2802_ | ~new_n2790_ | ~new_n2833_) & (new_n2802_ | ~new_n2790_ | ~new_n2826_) & ((~new_n2790_ & ~new_n2796_) | new_n2802_ | ~new_n2809_) & (~new_n2796_ | new_n2821_ | (new_n2790_ & new_n2833_)) & (new_n2833_ | ((~new_n2802_ | new_n2809_) & ~new_n2826_ & (new_n2790_ | new_n2796_))) & (new_n2815_ | (new_n2821_ & (new_n2790_ ? new_n2826_ : ~new_n2796_))) & ((new_n2802_ ^ new_n2809_) | ~new_n2826_ | ~new_n2833_ | ~new_n2815_ | ~new_n2821_ | new_n2790_ | ~new_n2796_) & (~new_n2802_ | ~new_n2790_ | ~new_n2821_ | ~new_n2826_ | ~new_n2833_ | ~new_n2796_ | new_n2815_) & (new_n2802_ | ~new_n2809_ | ~new_n2833_ | new_n2790_ | new_n2796_ | ~new_n2815_ | new_n2826_ | new_n2821_) & (~new_n2826_ | ~new_n2821_ | ~new_n2833_ | new_n2790_ | new_n2796_ | new_n2815_ | new_n2802_ | ~new_n2809_) & (~new_n2790_ | ~new_n2821_ | ~new_n2802_ | ~new_n2809_ | new_n2826_ | ~new_n2815_ | new_n2833_);
  assign new_n3287_ = (~new_n2802_ | ~new_n2833_ | new_n2790_ | new_n2796_ | new_n2826_ | ~new_n2821_ | ~new_n2809_ | new_n2815_) & (~new_n2815_ | new_n2826_ | new_n2821_ | ~new_n2796_ | new_n2809_ | ~new_n2790_ | ~new_n2833_) & (new_n2826_ | ~new_n2821_ | ~new_n2833_ | new_n2790_ | new_n2796_ | new_n2815_ | new_n2802_ | ~new_n2809_) & (new_n2826_ | ~new_n2802_ | ~new_n2809_ | ~new_n2815_ | ~new_n2821_ | new_n2790_ | ~new_n2796_);
  assign new_n3288_ = ((new_n2925_ & ~P3_INSTADDRPOINTER_REG_15__SCAN_IN) | (~new_n2925_ & P3_INSTADDRPOINTER_REG_15__SCAN_IN) | ((new_n2925_ | ~P3_INSTADDRPOINTER_REG_14__SCAN_IN) & (new_n2931_ | (new_n2925_ & ~P3_INSTADDRPOINTER_REG_14__SCAN_IN)))) & new_n3289_ & ((new_n2925_ ^ ~P3_INSTADDRPOINTER_REG_15__SCAN_IN) | (~new_n2925_ & P3_INSTADDRPOINTER_REG_14__SCAN_IN) | (~new_n2931_ & (~new_n2925_ | P3_INSTADDRPOINTER_REG_14__SCAN_IN)));
  assign new_n3289_ = ~new_n2906_ & ~new_n2802_ & new_n2950_ & ((new_n2927_ & new_n2939_) | (new_n2928_ & new_n2945_));
  assign new_n3290_ = ((P3_INSTADDRPOINTER_REG_15__SCAN_IN & new_n3278_ & new_n2782_) | ~new_n3306_ | (~P3_INSTADDRPOINTER_REG_15__SCAN_IN & (~new_n3278_ | ~new_n2782_))) & new_n3292_ & ((new_n3291_ & P3_INSTADDRPOINTER_REG_15__SCAN_IN) | ~new_n3307_ | (~new_n3291_ & ~P3_INSTADDRPOINTER_REG_15__SCAN_IN));
  assign new_n3291_ = new_n2782_ & new_n2924_ & (new_n2913_ | ~new_n2922_);
  assign new_n3292_ = (new_n3296_ | (~P3_PHYADDRPOINTER_REG_15__SCAN_IN ^ (P3_PHYADDRPOINTER_REG_1__SCAN_IN & new_n3299_ & P3_PHYADDRPOINTER_REG_14__SCAN_IN))) & ~new_n3304_ & (~new_n3293_ | ~P3_PHYADDRPOINTER_REG_15__SCAN_IN) & (new_n3293_ | ~new_n3305_ | (P3_PHYADDRPOINTER_REG_15__SCAN_IN & new_n3299_ & P3_PHYADDRPOINTER_REG_14__SCAN_IN) | (~P3_PHYADDRPOINTER_REG_15__SCAN_IN & (~new_n3299_ | ~P3_PHYADDRPOINTER_REG_14__SCAN_IN)));
  assign new_n3293_ = ~new_n3294_ & (~new_n2950_ | ((~new_n2927_ | ~new_n2939_) & (~new_n2928_ | ~new_n2945_)));
  assign new_n3294_ = new_n3283_ & ~new_n3295_;
  assign new_n3295_ = P3_STATE2_REG_2__SCAN_IN & P3_STATE2_REG_1__SCAN_IN;
  assign new_n3296_ = (~new_n3297_ | (~new_n3294_ & (~new_n2950_ | ((~new_n2927_ | ~new_n2939_) & (~new_n2928_ | ~new_n2945_))))) & (~new_n3298_ | (~new_n3294_ & (~new_n2950_ | ((~new_n2927_ | ~new_n2939_) & (~new_n2928_ | ~new_n2945_)))));
  assign new_n3297_ = P3_STATE2_REG_2__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN;
  assign new_n3298_ = P3_STATE2_REG_1__SCAN_IN & ~P3_STATEBS16_REG_SCAN_IN;
  assign new_n3299_ = P3_PHYADDRPOINTER_REG_13__SCAN_IN & new_n3300_ & P3_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign new_n3300_ = new_n3301_ & P3_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign new_n3301_ = new_n3302_ & new_n3303_;
  assign new_n3302_ = P3_PHYADDRPOINTER_REG_6__SCAN_IN & P3_PHYADDRPOINTER_REG_5__SCAN_IN & P3_PHYADDRPOINTER_REG_4__SCAN_IN & P3_PHYADDRPOINTER_REG_2__SCAN_IN & P3_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign new_n3303_ = P3_PHYADDRPOINTER_REG_10__SCAN_IN & P3_PHYADDRPOINTER_REG_9__SCAN_IN & P3_PHYADDRPOINTER_REG_7__SCAN_IN & P3_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign new_n3304_ = P3_REIP_REG_15__SCAN_IN & new_n3284_ & (new_n3294_ | (new_n2950_ & ((new_n2927_ & new_n2939_) | (new_n2928_ & new_n2945_))));
  assign new_n3305_ = P3_STATE2_REG_1__SCAN_IN & P3_STATEBS16_REG_SCAN_IN;
  assign new_n3306_ = new_n2802_ & new_n2950_ & ((new_n2927_ & new_n2939_) | (new_n2928_ & new_n2945_));
  assign new_n3307_ = new_n2906_ & ~new_n2802_ & new_n2950_ & ((new_n2927_ & new_n2939_) | (new_n2928_ & new_n2945_));
  assign new_n3308_ = (new_n1678_ | new_n1672_ | new_n1667_) & new_n2706_ & (new_n2667_ | new_n2684_ | (new_n1787_ & new_n1764_));
  assign new_n3309_ = ~P1_EBX_REG_4__SCAN_IN & ~P1_EBX_REG_1__SCAN_IN & ~P1_EBX_REG_19__SCAN_IN & ~P1_EBX_REG_12__SCAN_IN;
  assign new_n3310_ = (~new_n3311_ | P1_REQUESTPENDING_REG_SCAN_IN) & (new_n3311_ | ~new_n3314_) & (~new_n2690_ | ~new_n3313_) & (new_n2723_ | new_n3315_);
  assign new_n3311_ = (~new_n2118_ | (~new_n2631_ & new_n2632_)) & ~new_n2119_ & ~new_n2576_ & (new_n2510_ | ~new_n3312_);
  assign new_n3312_ = P1_STATE2_REG_1__SCAN_IN & P1_STATE2_REG_2__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN;
  assign new_n3313_ = ~new_n1982_ ^ (~new_n1981_ & (new_n1979_ | (~new_n1980_ & (new_n1383_ | (~new_n1386_ & ~new_n1387_)))));
  assign new_n3314_ = (~P1_STATE2_REG_0__SCAN_IN | (~new_n2510_ & P1_STATE2_REG_2__SCAN_IN & (~new_n2067_ | new_n2073_ | (new_n2567_ & P1_STATEBS16_REG_SCAN_IN)))) & (P1_STATE2_REG_2__SCAN_IN | P1_STATE2_REG_1__SCAN_IN) & (new_n2567_ | ~P1_STATE2_REG_0__SCAN_IN | new_n2067_ | ~new_n2073_);
  assign new_n3315_ = ~P2_EBX_REG_13__SCAN_IN & ~P2_EBX_REG_15__SCAN_IN & ~P2_EBX_REG_20__SCAN_IN & ~P2_EBX_REG_22__SCAN_IN & ~P2_EBX_REG_25__SCAN_IN & ~P2_EBX_REG_31__SCAN_IN;
  assign new_n3316_ = new_n3317_ & (new_n3050_ | ~new_n2505_ | ~new_n2513_) & (~new_n2584_ | (new_n2578_ & P1_INSTADDRPOINTER_REG_17__SCAN_IN) | (~new_n2578_ & ~P1_INSTADDRPOINTER_REG_17__SCAN_IN));
  assign new_n3317_ = (new_n3318_ | new_n2587_ | ~new_n2495_ | (~new_n2566_ & new_n2568_)) & (new_n3319_ | new_n2575_ | (new_n2495_ & (new_n2566_ | ~new_n2568_)));
  assign new_n3318_ = ((~P1_INSTADDRPOINTER_REG_20__SCAN_IN & (~P1_INSTADDRPOINTER_REG_0__SCAN_IN | ~new_n2583_ | ~P1_INSTADDRPOINTER_REG_17__SCAN_IN | ~P1_INSTADDRPOINTER_REG_16__SCAN_IN | ~P1_INSTADDRPOINTER_REG_15__SCAN_IN | ~new_n2579_ | ~P1_INSTADDRPOINTER_REG_14__SCAN_IN)) | (P1_INSTADDRPOINTER_REG_0__SCAN_IN & P1_INSTADDRPOINTER_REG_20__SCAN_IN & new_n2583_ & P1_INSTADDRPOINTER_REG_17__SCAN_IN & P1_INSTADDRPOINTER_REG_16__SCAN_IN & P1_INSTADDRPOINTER_REG_15__SCAN_IN & new_n2579_ & P1_INSTADDRPOINTER_REG_14__SCAN_IN)) & (~P1_INSTADDRPOINTER_REG_17__SCAN_IN | (P1_INSTADDRPOINTER_REG_16__SCAN_IN & P1_INSTADDRPOINTER_REG_15__SCAN_IN & P1_INSTADDRPOINTER_REG_14__SCAN_IN & new_n2579_ & P1_INSTADDRPOINTER_REG_0__SCAN_IN)) & (P1_INSTADDRPOINTER_REG_17__SCAN_IN | ~P1_INSTADDRPOINTER_REG_16__SCAN_IN | ~P1_INSTADDRPOINTER_REG_15__SCAN_IN | ~P1_INSTADDRPOINTER_REG_14__SCAN_IN | ~new_n2579_ | ~P1_INSTADDRPOINTER_REG_0__SCAN_IN);
  assign new_n3319_ = ~P1_INSTADDRPOINTER_REG_16__SCAN_IN & ~P1_INSTADDRPOINTER_REG_14__SCAN_IN & ~P1_INSTADDRPOINTER_REG_20__SCAN_IN & ~P1_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign new_n3320_ = ~new_n3321_ & ((new_n2986_ & ~new_n3148_) | new_n2067_ | ~new_n2073_ | new_n2630_ | ~P1_STATE2_REG_2__SCAN_IN);
  assign new_n3321_ = ((~P3_INSTADDRPOINTER_REG_11__SCAN_IN & (~new_n3278_ | ~P3_INSTADDRPOINTER_REG_10__SCAN_IN)) | ~new_n3306_ | (new_n3278_ & P3_INSTADDRPOINTER_REG_10__SCAN_IN & P3_INSTADDRPOINTER_REG_11__SCAN_IN)) & ~new_n3322_ & ~new_n3323_ & new_n3324_;
  assign new_n3322_ = (((~new_n2925_ | P3_INSTADDRPOINTER_REG_10__SCAN_IN) & (new_n2913_ | ~new_n2932_) & (~new_n2925_ | (P3_INSTADDRPOINTER_REG_8__SCAN_IN & P3_INSTADDRPOINTER_REG_9__SCAN_IN))) | (~new_n2925_ & P3_INSTADDRPOINTER_REG_9__SCAN_IN) | (~new_n2925_ & P3_INSTADDRPOINTER_REG_10__SCAN_IN) | (new_n2925_ ^ ~P3_INSTADDRPOINTER_REG_11__SCAN_IN)) & new_n3289_ & ((((new_n2925_ & ~P3_INSTADDRPOINTER_REG_10__SCAN_IN) | (~new_n2913_ & new_n2932_) | (new_n2925_ & (~P3_INSTADDRPOINTER_REG_8__SCAN_IN | ~P3_INSTADDRPOINTER_REG_9__SCAN_IN))) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_9__SCAN_IN) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_10__SCAN_IN)) | (new_n2925_ & ~P3_INSTADDRPOINTER_REG_11__SCAN_IN) | (~new_n2925_ & P3_INSTADDRPOINTER_REG_11__SCAN_IN));
  assign new_n3323_ = (P3_INSTADDRPOINTER_REG_11__SCAN_IN | (P3_INSTADDRPOINTER_REG_10__SCAN_IN & new_n2924_ & (new_n2913_ | ~new_n2922_))) & new_n3307_ & (~P3_INSTADDRPOINTER_REG_10__SCAN_IN | ~P3_INSTADDRPOINTER_REG_11__SCAN_IN | ~new_n2924_ | (~new_n2913_ & new_n2922_));
  assign new_n3324_ = (new_n3296_ | (~P3_PHYADDRPOINTER_REG_11__SCAN_IN ^ (new_n3301_ & P3_PHYADDRPOINTER_REG_1__SCAN_IN))) & (new_n3293_ | ~new_n3284_ | ~P3_REIP_REG_11__SCAN_IN) & (~new_n3293_ | ~P3_PHYADDRPOINTER_REG_11__SCAN_IN) & (new_n3293_ | ~new_n3305_ | (new_n3301_ & P3_PHYADDRPOINTER_REG_11__SCAN_IN) | (~new_n3301_ & ~P3_PHYADDRPOINTER_REG_11__SCAN_IN));
  assign new_n3325_ = new_n3326_ & ~new_n3329_ & (~new_n2586_ | (P1_INSTADDRPOINTER_REG_16__SCAN_IN & P1_INSTADDRPOINTER_REG_15__SCAN_IN & P1_INSTADDRPOINTER_REG_14__SCAN_IN & new_n2579_ & P1_INSTADDRPOINTER_REG_0__SCAN_IN) | (~P1_INSTADDRPOINTER_REG_16__SCAN_IN & (~P1_INSTADDRPOINTER_REG_15__SCAN_IN | ~P1_INSTADDRPOINTER_REG_14__SCAN_IN | ~new_n2579_ | ~P1_INSTADDRPOINTER_REG_0__SCAN_IN)));
  assign new_n3326_ = (new_n3328_ | ~new_n2493_ | ~new_n2495_ | (~new_n2566_ & new_n2568_)) & (~new_n3327_ | ~new_n2585_ | ~new_n2495_ | (~new_n2566_ & new_n2568_));
  assign new_n3327_ = P1_INSTADDRPOINTER_REG_16__SCAN_IN ^ (P1_INSTADDRPOINTER_REG_15__SCAN_IN & new_n2579_ & P1_INSTADDRPOINTER_REG_14__SCAN_IN);
  assign new_n3328_ = (~new_n2593_ ^ P1_INSTADDRPOINTER_REG_14__SCAN_IN) & (~P1_INSTADDRPOINTER_REG_16__SCAN_IN ^ (P1_INSTADDRPOINTER_REG_15__SCAN_IN & new_n2593_ & P1_INSTADDRPOINTER_REG_14__SCAN_IN));
  assign new_n3329_ = ~new_n3330_ & new_n3333_ & ((~P3_INSTADDRPOINTER_REG_7__SCAN_IN & (~new_n2904_ ^ (~new_n2865_ ^ ~new_n2906_))) | ~new_n3306_ | ((new_n2904_ | (new_n2865_ & ~new_n2906_) | (~new_n2865_ & new_n2906_)) & P3_INSTADDRPOINTER_REG_7__SCAN_IN & (~new_n2904_ | (new_n2865_ ^ ~new_n2906_))));
  assign new_n3330_ = (~new_n3331_ | (~P3_INSTADDRPOINTER_REG_7__SCAN_IN & (new_n2923_ ^ new_n2906_)) | (P3_INSTADDRPOINTER_REG_7__SCAN_IN & (new_n2923_ | ~new_n2906_) & (~new_n2923_ | new_n2906_))) & new_n3332_ & (new_n3331_ | (~P3_INSTADDRPOINTER_REG_7__SCAN_IN ^ (new_n2923_ ^ new_n2906_)));
  assign new_n3331_ = ~new_n2915_ & (~new_n2921_ | (~new_n2916_ & (new_n2918_ | ~new_n2920_) & (new_n2917_ | P3_INSTADDRPOINTER_REG_4__SCAN_IN)));
  assign new_n3332_ = ~new_n2802_ & new_n2950_ & ((new_n2927_ & new_n2939_) | (new_n2928_ & new_n2945_));
  assign new_n3333_ = (new_n3296_ | (~new_n3334_ & ~P3_PHYADDRPOINTER_REG_7__SCAN_IN) | (new_n3334_ & P3_PHYADDRPOINTER_REG_7__SCAN_IN)) & (new_n3293_ | ~new_n3305_ | (new_n3302_ & P3_PHYADDRPOINTER_REG_7__SCAN_IN) | (~new_n3302_ & ~P3_PHYADDRPOINTER_REG_7__SCAN_IN)) & (~new_n3293_ | ~P3_PHYADDRPOINTER_REG_7__SCAN_IN) & (~P3_REIP_REG_7__SCAN_IN | new_n3293_ | ~new_n3284_);
  assign new_n3334_ = P3_PHYADDRPOINTER_REG_6__SCAN_IN & P3_PHYADDRPOINTER_REG_1__SCAN_IN & P3_PHYADDRPOINTER_REG_5__SCAN_IN & P3_PHYADDRPOINTER_REG_4__SCAN_IN & P3_PHYADDRPOINTER_REG_2__SCAN_IN & P3_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign new_n3335_ = new_n3336_ & (~new_n2630_ | new_n3339_) & (~new_n2505_ | ~new_n2513_ | (new_n2954_ ? ~BUF1_REG_0__SCAN_IN : ~DATAI_0_));
  assign new_n3336_ = (~new_n3337_ | new_n2587_ | ~new_n2495_ | (~new_n2566_ & new_n2568_)) & (~new_n3338_ | new_n2572_ | ~new_n2495_ | (~new_n2566_ & new_n2568_));
  assign new_n3337_ = P1_INSTADDRPOINTER_REG_14__SCAN_IN ^ (new_n2579_ & P1_INSTADDRPOINTER_REG_0__SCAN_IN);
  assign new_n3338_ = new_n2454_ ^ (~new_n2469_ & new_n2468_ & new_n2467_ & new_n2457_ & new_n2463_);
  assign new_n3339_ = ~P1_REIP_REG_1__SCAN_IN & ~P1_REIP_REG_23__SCAN_IN & ~P1_REIP_REG_22__SCAN_IN;
  assign new_n3340_ = new_n3341_ & ~new_n3348_ & (new_n3156_ | ~new_n2505_ | ~new_n2291_) & new_n3350_ & ~new_n3354_ & (new_n3123_ | ~new_n2505_ | ~new_n2291_);
  assign new_n3341_ = ~new_n3342_ & ((~P1_REIP_REG_4__SCAN_IN & ~P1_REIP_REG_19__SCAN_IN & ~P1_REIP_REG_12__SCAN_IN) | ~new_n2633_ | (new_n2118_ & (new_n2631_ | ~new_n2632_)));
  assign new_n3342_ = (~new_n3347_ | ~new_n3346_ | (~new_n3343_ & ~new_n3344_ & ~new_n3345_ & (new_n2913_ | ~new_n2932_))) & new_n3289_ & (new_n3347_ | (new_n3346_ & (new_n3343_ | new_n3344_ | new_n3345_ | (~new_n2913_ & new_n2932_))));
  assign new_n3343_ = new_n2925_ & ~P3_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign new_n3344_ = new_n2925_ & ~P3_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign new_n3345_ = new_n2925_ & ~new_n2784_;
  assign new_n3346_ = (new_n2925_ | ~P3_INSTADDRPOINTER_REG_11__SCAN_IN) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_9__SCAN_IN) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  assign new_n3347_ = new_n2925_ ^ P3_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign new_n3348_ = new_n2509_ & ((P1_EAX_REG_9__SCAN_IN & new_n3349_ & new_n2067_) | (new_n3349_ & ~new_n2067_ & (new_n2954_ | DATAI_9_) & (~new_n2954_ | BUF1_REG_9__SCAN_IN)));
  assign new_n3349_ = new_n2495_ & ~new_n2073_ & (new_n2478_ | new_n2482_) & (~new_n2510_ | (new_n2067_ & ~new_n2073_));
  assign new_n3350_ = (~new_n2991_ | (~new_n3013_ & ~new_n3351_)) & (~new_n3353_ | (~new_n3056_ & ~new_n3352_));
  assign new_n3351_ = ~new_n2085_ & P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN & (new_n2997_ | (P1_STATE2_REG_3__SCAN_IN & (new_n2478_ | new_n2482_)));
  assign new_n3352_ = ~new_n2073_ & P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN & (new_n2997_ | (P1_STATE2_REG_3__SCAN_IN & (new_n2478_ | new_n2482_)));
  assign new_n3353_ = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n3354_ = new_n3100_ & ((~new_n2067_ & P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN & (new_n2997_ | (~new_n2477_ & P1_STATE2_REG_3__SCAN_IN))) | (~new_n2079_ & P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN & (new_n2997_ | (~new_n2477_ & P1_STATE2_REG_3__SCAN_IN))));
  assign new_n3355_ = new_n3356_ & ((~P1_EBX_REG_23__SCAN_IN & ~P1_EBX_REG_22__SCAN_IN) | (~new_n2641_ & ~new_n2642_));
  assign new_n3356_ = (~new_n2448_ | ~new_n3359_) & ((new_n3358_ & P3_INSTADDRPOINTER_REG_12__SCAN_IN) | ~new_n3306_ | (~new_n3358_ & ~P3_INSTADDRPOINTER_REG_12__SCAN_IN)) & ((~P3_INSTADDRPOINTER_REG_21__SCAN_IN & (~new_n3357_ | ~new_n2787_)) | ~new_n3306_ | (new_n3357_ & new_n2787_ & P3_INSTADDRPOINTER_REG_21__SCAN_IN));
  assign new_n3357_ = new_n2781_ & ((P3_INSTADDRPOINTER_REG_7__SCAN_IN & (~new_n2904_ | (new_n2865_ ^ ~new_n2906_))) | (~new_n2904_ & (~new_n2865_ | new_n2906_) & (new_n2865_ | ~new_n2906_)) | (P3_INSTADDRPOINTER_REG_8__SCAN_IN & new_n2865_ & ~new_n2906_)) & P3_INSTADDRPOINTER_REG_9__SCAN_IN & (P3_INSTADDRPOINTER_REG_8__SCAN_IN | (new_n2865_ & ~new_n2906_));
  assign new_n3358_ = P3_INSTADDRPOINTER_REG_10__SCAN_IN & P3_INSTADDRPOINTER_REG_11__SCAN_IN & ((P3_INSTADDRPOINTER_REG_7__SCAN_IN & (~new_n2904_ | (new_n2865_ ^ ~new_n2906_))) | (P3_INSTADDRPOINTER_REG_8__SCAN_IN & new_n2865_ & ~new_n2906_) | (~new_n2904_ & (~new_n2865_ | new_n2906_) & (new_n2865_ | ~new_n2906_))) & P3_INSTADDRPOINTER_REG_9__SCAN_IN & (P3_INSTADDRPOINTER_REG_8__SCAN_IN | (new_n2865_ & ~new_n2906_));
  assign new_n3359_ = ~new_n3360_ & (new_n2606_ | (new_n2605_ & ~new_n2073_ & (new_n2478_ | new_n2482_)));
  assign new_n3360_ = (~P1_STATE2_REG_2__SCAN_IN | P1_STATE2_REG_0__SCAN_IN) & (P1_STATEBS16_REG_SCAN_IN | ~P1_STATE2_REG_1__SCAN_IN);
  assign new_n3361_ = (~new_n3199_ | ~new_n3211_) & (~new_n3082_ | (~new_n3189_ & ~new_n3244_));
  assign new_n3362_ = (new_n3363_ | (new_n3364_ & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_2__SCAN_IN) & new_n2966_ & ((~P2_STATE2_REG_3__SCAN_IN & (new_n1810_ | ~P2_STATE2_REG_2__SCAN_IN)) | (new_n3364_ & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN));
  assign new_n3363_ = P2_STATEBS16_REG_SCAN_IN & new_n1666_ & (~new_n1664_ | (new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_))) & (new_n1664_ | ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ ^ (~new_n1409_ ^ new_n1421_));
  assign new_n3364_ = P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3365_ = new_n3366_ & (~new_n2683_ | new_n1335_ | (~new_n1419_ & (new_n1662_ | new_n1420_)) | (new_n1419_ & ~new_n1662_ & ~new_n1420_));
  assign new_n3366_ = (~new_n3070_ | new_n1670_ | ~new_n1666_ | (new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) | (~new_n1412_ ^ (new_n1409_ ^ ~new_n1421_))) & (~new_n3195_ | new_n1670_ | new_n1666_ | (new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) | (~new_n1412_ ^ (new_n1409_ ^ ~new_n1421_)));
  assign new_n3367_ = new_n3383_ & new_n3377_ & ~new_n3368_ & ((new_n1657_ & new_n2665_) | ~new_n3372_ | ~new_n3375_);
  assign new_n3368_ = new_n3071_ & ((P2_STATE2_REG_2__SCAN_IN & (new_n1808_ | new_n3370_)) | ((~new_n3369_ | ~P2_STATEBS16_REG_SCAN_IN) & new_n3371_ & ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN));
  assign new_n3369_ = new_n1666_ & (~new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ ^ (~new_n1409_ ^ new_n1421_));
  assign new_n3370_ = P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3371_ = P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3372_ = new_n3373_ & (new_n2723_ | ~P2_EBX_REG_10__SCAN_IN) & (~new_n2756_ | (P2_PHYADDRPOINTER_REG_10__SCAN_IN & new_n2019_ & P2_PHYADDRPOINTER_REG_9__SCAN_IN) | (~P2_PHYADDRPOINTER_REG_10__SCAN_IN & (~new_n2019_ | ~P2_PHYADDRPOINTER_REG_9__SCAN_IN)));
  assign new_n3373_ = (~new_n2757_ | (new_n1914_ & new_n1915_) | (~new_n1914_ & ~new_n1915_)) & (~P2_PHYADDRPOINTER_REG_10__SCAN_IN | new_n2724_ | ~P2_STATE2_REG_3__SCAN_IN) & (new_n2724_ | ~new_n3374_) & (~new_n2724_ | ~P2_REIP_REG_10__SCAN_IN);
  assign new_n3374_ = new_n2970_ & ~P2_STATE2_REG_1__SCAN_IN;
  assign new_n3375_ = ~new_n3376_ & (~new_n2726_ | (~new_n2747_ & (~new_n2738_ | new_n2748_)) | (new_n2747_ & new_n2738_ & ~new_n2748_));
  assign new_n3376_ = (~new_n1987_ | (~new_n1986_ & ~new_n1985_ & new_n1978_ & ~new_n1984_)) & new_n2691_ & (new_n1987_ | new_n1986_ | new_n1985_ | ~new_n1978_ | new_n1984_);
  assign new_n3377_ = (new_n3379_ | ~new_n3166_) & ((~new_n3054_ & ~new_n3229_) | ~new_n3378_ | ~new_n2994_);
  assign new_n3378_ = (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ | (new_n2148_ & new_n2200_) | (~new_n2148_ & ~new_n2200_)) & (~new_n2154_ | (new_n2148_ ^ new_n2200_));
  assign new_n3379_ = ~new_n3380_ & (~new_n3382_ | (P2_STATEBS16_REG_SCAN_IN & new_n1666_ & (~new_n1664_ | (new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_))) & (new_n1664_ | ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ ^ (~new_n1409_ ^ new_n1421_))));
  assign new_n3380_ = P2_STATE2_REG_2__SCAN_IN & (new_n3381_ | (new_n1413_ & new_n1803_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_)) & (new_n1387_ ^ (~new_n1383_ & ~new_n1386_))));
  assign new_n3381_ = new_n3364_ & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n3382_ = new_n2970_ & new_n3364_ & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n3383_ = (~new_n3103_ | ~new_n3124_) & (~new_n3030_ | new_n3384_) & ~new_n3385_ & (~new_n3266_ | ~new_n3012_);
  assign new_n3384_ = ~new_n3165_ & (~new_n2996_ | (~new_n2954_ & ~DATAI_20_) | (new_n2954_ & ~BUF1_REG_20__SCAN_IN));
  assign new_n3385_ = ~new_n2630_ & ~new_n3386_ & (~new_n2287_ ^ (new_n2285_ ^ (~new_n2284_ | ~new_n2237_)));
  assign new_n3386_ = (new_n2644_ | ~P1_STATE2_REG_1__SCAN_IN) & (~P1_STATE2_REG_2__SCAN_IN | ~new_n2067_ | ~new_n2073_);
  assign new_n3387_ = ~new_n3396_ & (new_n3389_ | ~P2_INSTQUEUE_REG_3__4__SCAN_IN) & (~new_n3397_ | new_n3398_) & (~new_n3391_ | (~new_n3388_ & P2_INSTQUEUE_REG_5__4__SCAN_IN));
  assign new_n3388_ = ~new_n3233_ & new_n3235_;
  assign new_n3389_ = new_n3390_ & (new_n3371_ | (~new_n2969_ & (new_n3369_ | ~new_n2968_)));
  assign new_n3390_ = new_n2966_ & (new_n3370_ | (~P2_STATE2_REG_3__SCAN_IN & (new_n1808_ | ~P2_STATE2_REG_2__SCAN_IN)));
  assign new_n3391_ = (new_n3392_ | ~new_n3071_) & new_n3394_ & (~new_n3393_ | ~new_n3070_);
  assign new_n3392_ = ~new_n3238_ & (~new_n3239_ | (new_n3234_ & (~new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_))));
  assign new_n3393_ = new_n3242_ & (~new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_));
  assign new_n3394_ = ~new_n3395_ & (~new_n3069_ | ~new_n2963_ | (new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) | (~new_n1412_ & (~new_n1409_ | new_n1421_) & (new_n1409_ | ~new_n1421_)) | (new_n1412_ & (~new_n1409_ ^ ~new_n1421_)));
  assign new_n3395_ = new_n3236_ & ~new_n1350_ & new_n2966_ & P2_STATE2_REG_3__SCAN_IN;
  assign new_n3396_ = new_n2757_ & ((new_n1944_ ^ (new_n1942_ & (~new_n1330_ | ~P2_EBX_REG_19__SCAN_IN))) | (new_n1948_ ^ ((~new_n1330_ | ~P2_EBX_REG_21__SCAN_IN) & new_n1944_ & new_n1942_ & (~new_n1330_ | ~P2_EBX_REG_19__SCAN_IN))));
  assign new_n3397_ = ~new_n2994_ & new_n2284_ & (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & (new_n2154_ ^ (new_n2148_ ^ new_n2200_));
  assign new_n3398_ = ~new_n3104_ & ~new_n3165_;
  assign new_n3399_ = new_n3400_ & new_n3409_ & new_n4080_ & new_n3410_ & new_n4071_ & new_n3419_ & new_n3431_ & new_n4042_;
  assign new_n3400_ = (~new_n3402_ | ~new_n2691_) & (~new_n2639_ | new_n3406_) & ~new_n3403_ & (~new_n3401_ | (~new_n2659_ & new_n3404_));
  assign new_n3401_ = new_n2476_ & new_n2053_;
  assign new_n3402_ = ~new_n1991_ ^ (new_n1988_ & ~new_n1987_ & ~new_n1986_ & ~new_n1985_ & new_n1978_ & ~new_n1984_);
  assign new_n3403_ = (new_n2517_ | new_n2659_) & P1_EBX_REG_31__SCAN_IN & ~new_n2634_ & ~new_n2630_ & new_n2494_ & P1_STATE2_REG_2__SCAN_IN;
  assign new_n3404_ = (~new_n2453_ ^ new_n2473_) & (new_n3405_ ^ (new_n2453_ & new_n2473_));
  assign new_n3405_ = new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_20__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_20__SCAN_IN));
  assign new_n3406_ = new_n3408_ & ((~P1_REIP_REG_23__SCAN_IN & ~P1_REIP_REG_22__SCAN_IN & ((~new_n3407_ & ~P1_REIP_REG_19__SCAN_IN) | ((~P1_REIP_REG_21__SCAN_IN | ~P1_REIP_REG_20__SCAN_IN) & new_n3407_ & P1_REIP_REG_19__SCAN_IN))) | (new_n3407_ & P1_REIP_REG_19__SCAN_IN & P1_REIP_REG_23__SCAN_IN & P1_REIP_REG_22__SCAN_IN & P1_REIP_REG_21__SCAN_IN & P1_REIP_REG_20__SCAN_IN));
  assign new_n3407_ = P1_REIP_REG_18__SCAN_IN & P1_REIP_REG_15__SCAN_IN & P1_REIP_REG_17__SCAN_IN & P1_REIP_REG_16__SCAN_IN & P1_REIP_REG_14__SCAN_IN & new_n2646_ & P1_REIP_REG_13__SCAN_IN & P1_REIP_REG_12__SCAN_IN;
  assign new_n3408_ = (new_n2646_ | ~P1_REIP_REG_12__SCAN_IN) & (~new_n2646_ | P1_REIP_REG_12__SCAN_IN) & (P1_REIP_REG_4__SCAN_IN | ~P1_REIP_REG_3__SCAN_IN | ~P1_REIP_REG_2__SCAN_IN) & P1_REIP_REG_1__SCAN_IN & (~P1_REIP_REG_4__SCAN_IN | (P1_REIP_REG_3__SCAN_IN & P1_REIP_REG_2__SCAN_IN));
  assign new_n3409_ = (~new_n1657_ | ~new_n2678_) & (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | new_n3003_ | (new_n3151_ & (~new_n3147_ | (~new_n3130_ & new_n3138_))));
  assign new_n3410_ = new_n3418_ & ~new_n3411_ & (~new_n3058_ | ~new_n2968_ | ~new_n2981_);
  assign new_n3411_ = new_n2726_ & ((new_n3412_ & ~new_n3413_) | (~new_n3412_ & new_n3417_) | ~new_n3415_ | (new_n2733_ ^ new_n2755_));
  assign new_n3412_ = (~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN) & (P2_STATE2_REG_0__SCAN_IN | (P2_PHYADDRPOINTER_REG_24__SCAN_IN & new_n2730_ & P2_PHYADDRPOINTER_REG_23__SCAN_IN) | (~P2_PHYADDRPOINTER_REG_24__SCAN_IN & (~new_n2730_ | ~P2_PHYADDRPOINTER_REG_23__SCAN_IN))) & new_n2733_ & new_n2755_ & (~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN) & (P2_STATE2_REG_0__SCAN_IN | (~new_n2730_ & ~P2_PHYADDRPOINTER_REG_23__SCAN_IN) | (new_n2730_ & P2_PHYADDRPOINTER_REG_23__SCAN_IN));
  assign new_n3413_ = (new_n3414_ | P2_STATE2_REG_0__SCAN_IN) & (~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_25__SCAN_IN) & (~P2_STATE2_REG_0__SCAN_IN | P2_INSTADDRPOINTER_REG_26__SCAN_IN | P2_INSTADDRPOINTER_REG_27__SCAN_IN | P2_INSTADDRPOINTER_REG_28__SCAN_IN | P2_INSTADDRPOINTER_REG_29__SCAN_IN | P2_INSTADDRPOINTER_REG_30__SCAN_IN);
  assign new_n3414_ = (~P2_PHYADDRPOINTER_REG_30__SCAN_IN | ~P2_PHYADDRPOINTER_REG_29__SCAN_IN | ~P2_PHYADDRPOINTER_REG_28__SCAN_IN | ~P2_PHYADDRPOINTER_REG_26__SCAN_IN | ~P2_PHYADDRPOINTER_REG_27__SCAN_IN | ~new_n2016_ | ~P2_PHYADDRPOINTER_REG_25__SCAN_IN) & (~new_n2016_ ^ P2_PHYADDRPOINTER_REG_25__SCAN_IN) & ((P2_PHYADDRPOINTER_REG_26__SCAN_IN & P2_PHYADDRPOINTER_REG_27__SCAN_IN & new_n2016_ & P2_PHYADDRPOINTER_REG_25__SCAN_IN) | new_n2016_ | P2_PHYADDRPOINTER_REG_25__SCAN_IN | P2_PHYADDRPOINTER_REG_26__SCAN_IN | P2_PHYADDRPOINTER_REG_27__SCAN_IN | P2_PHYADDRPOINTER_REG_30__SCAN_IN | P2_PHYADDRPOINTER_REG_28__SCAN_IN | P2_PHYADDRPOINTER_REG_29__SCAN_IN);
  assign new_n3415_ = new_n3416_ & (~new_n2734_ ^ (new_n2764_ & new_n2753_));
  assign new_n3416_ = ((new_n2737_ | new_n2750_) ^ (new_n2746_ & ~new_n2744_ & ~new_n2749_ & new_n2747_ & new_n2738_ & ~new_n2748_)) & (new_n2744_ ^ (~new_n2749_ & new_n2747_ & new_n2738_ & ~new_n2748_));
  assign new_n3417_ = P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_25__SCAN_IN : (~new_n2016_ ^ P2_PHYADDRPOINTER_REG_25__SCAN_IN);
  assign new_n3418_ = (~new_n2968_ | new_n3194_ | ~new_n3059_ | (new_n1664_ & (~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_))) | (~new_n1664_ & ((new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_)))) | (~new_n1412_ & (new_n1409_ | ~new_n1421_) & (~new_n1409_ | new_n1421_)) | (new_n1412_ & (new_n1409_ ^ new_n1421_))) & (~new_n2968_ | ~new_n3210_ | ~new_n3059_ | (new_n1664_ & (~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_))) | (~new_n1664_ & ((new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_)))) | (~new_n1412_ ^ (~new_n1409_ ^ new_n1421_)));
  assign new_n3419_ = ~new_n3420_ & ~new_n3421_ & ~new_n3428_ & ~new_n3422_ & ~new_n3429_ & ~new_n3427_ & (~new_n3423_ | new_n3430_);
  assign new_n3420_ = new_n2757_ & (((new_n1925_ | ~new_n1330_ | ~P2_EBX_REG_13__SCAN_IN) & ~new_n1907_ & (~new_n1925_ | (new_n1330_ & P2_EBX_REG_13__SCAN_IN))) | ((~new_n1330_ | ~P2_EBX_REG_15__SCAN_IN | (new_n1925_ & (~new_n1330_ | ~P2_EBX_REG_13__SCAN_IN) & ~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_14__SCAN_IN))) & ~new_n1907_ & ((new_n1330_ & P2_EBX_REG_15__SCAN_IN) | ~new_n1925_ | (new_n1330_ & P2_EBX_REG_13__SCAN_IN) | new_n1907_ | (new_n1330_ & P2_EBX_REG_14__SCAN_IN))));
  assign new_n3421_ = P1_PHYADDRPOINTER_REG_1__SCAN_IN & ~new_n2630_ & P1_STATE2_REG_3__SCAN_IN;
  assign new_n3422_ = new_n2589_ & (P1_REIP_REG_16__SCAN_IN | P1_REIP_REG_20__SCAN_IN | P1_REIP_REG_17__SCAN_IN);
  assign new_n3423_ = ((~new_n2931_ & (~new_n2925_ | P3_INSTADDRPOINTER_REG_14__SCAN_IN) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_14__SCAN_IN)) | ~new_n3289_ | (new_n2931_ & (~new_n2925_ ^ ~P3_INSTADDRPOINTER_REG_14__SCAN_IN))) & new_n3426_ & (new_n3291_ | ~new_n3307_ | (~new_n3424_ & ~P3_INSTADDRPOINTER_REG_14__SCAN_IN));
  assign new_n3424_ = P3_INSTADDRPOINTER_REG_13__SCAN_IN & new_n3425_ & P3_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign new_n3425_ = P3_INSTADDRPOINTER_REG_10__SCAN_IN & P3_INSTADDRPOINTER_REG_11__SCAN_IN & new_n2924_ & (new_n2913_ | ~new_n2922_);
  assign new_n3426_ = (new_n3293_ | ~new_n3284_ | ~P3_REIP_REG_14__SCAN_IN) & (~new_n3293_ | ~P3_PHYADDRPOINTER_REG_14__SCAN_IN) & (new_n3293_ | ~new_n3305_ | (new_n3299_ & P3_PHYADDRPOINTER_REG_14__SCAN_IN) | (~new_n3299_ & ~P3_PHYADDRPOINTER_REG_14__SCAN_IN)) & (new_n3296_ | (~P3_PHYADDRPOINTER_REG_14__SCAN_IN & (~new_n3299_ | ~P3_PHYADDRPOINTER_REG_1__SCAN_IN)) | (P3_PHYADDRPOINTER_REG_1__SCAN_IN & new_n3299_ & P3_PHYADDRPOINTER_REG_14__SCAN_IN));
  assign new_n3427_ = new_n2565_ & ~new_n2572_ & (new_n2699_ | (~new_n3405_ ^ (new_n2453_ & new_n2473_)));
  assign new_n3428_ = (~new_n2509_ | ((~P1_EAX_REG_13__SCAN_IN | ~new_n3349_ | ~new_n2067_) & (~new_n3349_ | new_n2067_ | (~new_n2954_ & ~DATAI_13_) | (new_n2954_ & ~BUF1_REG_13__SCAN_IN)))) & (~P1_LWORD_REG_13__SCAN_IN | (new_n3349_ & new_n2509_));
  assign new_n3429_ = (~P1_UWORD_REG_1__SCAN_IN | (new_n3349_ & new_n2509_)) & (~new_n2509_ | ((~P1_EAX_REG_17__SCAN_IN | ~new_n3349_ | ~new_n2067_) & (~new_n3349_ | new_n2067_ | (new_n2954_ ? ~BUF1_REG_1__SCAN_IN : ~DATAI_1_))));
  assign new_n3430_ = new_n3306_ & (~new_n3278_ | ~new_n2782_) & (P3_INSTADDRPOINTER_REG_14__SCAN_IN | (new_n3358_ & new_n2934_));
  assign new_n3431_ = new_n4024_ & new_n3432_ & new_n3465_ & new_n3507_ & new_n3531_ & new_n3539_ & new_n3545_ & new_n3987_;
  assign new_n3432_ = new_n3436_ & ~new_n3433_ & ~new_n3434_ & ~new_n3438_ & ~new_n3441_ & ~new_n3442_ & (~new_n3176_ | new_n3464_);
  assign new_n3433_ = new_n3359_ & (new_n2246_ | new_n2259_);
  assign new_n3434_ = (P1_INSTQUEUE_REG_2__1__SCAN_IN | P1_INSTQUEUE_REG_2__6__SCAN_IN) & (~new_n3435_ | P1_STATE2_REG_0__SCAN_IN | (~new_n2997_ & (new_n2477_ | ~P1_STATE2_REG_3__SCAN_IN)));
  assign new_n3435_ = (~P1_STATE2_REG_2__SCAN_IN | (new_n2992_ & (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN))) & (~P1_STATE2_REG_3__SCAN_IN | (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & new_n2992_ & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN));
  assign new_n3436_ = (~new_n3359_ | ~new_n2438_) & (~new_n3437_ | ~P1_STATE2_REG_3__SCAN_IN | P1_STATE2_REG_0__SCAN_IN | (~new_n2997_ & (new_n2477_ | ~P1_STATE2_REG_3__SCAN_IN)));
  assign new_n3437_ = new_n3046_ & (~new_n2053_ | ~new_n2073_ | ~new_n2091_);
  assign new_n3438_ = (P2_UWORD_REG_4__SCAN_IN | P2_LWORD_REG_10__SCAN_IN | P2_LWORD_REG_7__SCAN_IN) & ~P2_STATE2_REG_0__SCAN_IN & (new_n3439_ | (P2_STATE2_REG_2__SCAN_IN & P2_STATE2_REG_1__SCAN_IN));
  assign new_n3439_ = new_n2670_ & (new_n3440_ | (new_n1791_ & new_n2667_ & ~new_n1762_ & (new_n1768_ | ~new_n1781_)));
  assign new_n3440_ = new_n1322_ & new_n1340_ & new_n1792_ & new_n1788_ & new_n1330_ & new_n1377_ & new_n1350_ & new_n1356_;
  assign new_n3441_ = ~new_n1317_ & new_n1759_ & ~new_n1335_ & (new_n2976_ ? BUF1_REG_22__SCAN_IN : BUF2_REG_22__SCAN_IN);
  assign new_n3442_ = new_n3443_ & (((~P3_PHYADDRPOINTER_REG_30__SCAN_IN | ~P3_PHYADDRPOINTER_REG_28__SCAN_IN | ~P3_PHYADDRPOINTER_REG_29__SCAN_IN | ~new_n3462_ | ~P3_PHYADDRPOINTER_REG_27__SCAN_IN) & (P3_PHYADDRPOINTER_REG_30__SCAN_IN | (P3_PHYADDRPOINTER_REG_28__SCAN_IN & P3_PHYADDRPOINTER_REG_29__SCAN_IN & new_n3462_ & P3_PHYADDRPOINTER_REG_27__SCAN_IN)) & new_n3463_ & (new_n3462_ ^ ~P3_PHYADDRPOINTER_REG_27__SCAN_IN) & ((new_n3462_ & P3_PHYADDRPOINTER_REG_27__SCAN_IN) ? (P3_PHYADDRPOINTER_REG_28__SCAN_IN & P3_PHYADDRPOINTER_REG_29__SCAN_IN) : (~P3_PHYADDRPOINTER_REG_28__SCAN_IN & ~P3_PHYADDRPOINTER_REG_29__SCAN_IN))) | ~new_n3453_ | ((~P3_PHYADDRPOINTER_REG_30__SCAN_IN ^ (P3_PHYADDRPOINTER_REG_28__SCAN_IN & P3_PHYADDRPOINTER_REG_29__SCAN_IN & new_n3462_ & P3_PHYADDRPOINTER_REG_27__SCAN_IN)) & (~new_n3463_ | (~new_n3462_ ^ ~P3_PHYADDRPOINTER_REG_27__SCAN_IN) | ((new_n3462_ & P3_PHYADDRPOINTER_REG_27__SCAN_IN) ? (~P3_PHYADDRPOINTER_REG_28__SCAN_IN | ~P3_PHYADDRPOINTER_REG_29__SCAN_IN) : (P3_PHYADDRPOINTER_REG_28__SCAN_IN | P3_PHYADDRPOINTER_REG_29__SCAN_IN)))));
  assign new_n3443_ = new_n3449_ & ~new_n3444_ & P3_STATE2_REG_1__SCAN_IN;
  assign new_n3444_ = new_n3448_ & (~new_n3445_ | new_n3447_);
  assign new_n3445_ = new_n3446_ & new_n2950_;
  assign new_n3446_ = ((~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) | (~new_n2940_ & (~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN))) & (~new_n2944_ | (new_n2940_ & (P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) & (~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)) | (~new_n2940_ & (P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ^ P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN)));
  assign new_n3447_ = (new_n2826_ | ~new_n2821_ | ~new_n2833_ | new_n2790_ | new_n2796_ | new_n2815_ | new_n2802_ | ~new_n2809_) & (~new_n2802_ | ~new_n2833_ | new_n2790_ | new_n2796_ | new_n2826_ | ~new_n2821_ | ~new_n2809_ | new_n2815_) & (~new_n2815_ | new_n2826_ | new_n2821_ | ~new_n2796_ | new_n2809_ | ~new_n2790_ | ~new_n2833_);
  assign new_n3448_ = (P3_STATE2_REG_2__SCAN_IN | P3_STATE2_REG_1__SCAN_IN | ~P3_STATE2_REG_3__SCAN_IN | ~P3_STATE2_REG_0__SCAN_IN) & (P3_STATE2_REG_2__SCAN_IN | P3_STATE2_REG_1__SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_0__SCAN_IN) & (~P3_STATE2_REG_1__SCAN_IN | P3_STATEBS16_REG_SCAN_IN | P3_STATE2_REG_2__SCAN_IN | P3_STATE2_REG_0__SCAN_IN);
  assign new_n3449_ = ~P3_PHYADDRPOINTER_REG_31__SCAN_IN ^ (~P3_PHYADDRPOINTER_REG_30__SCAN_IN | ~P3_PHYADDRPOINTER_REG_28__SCAN_IN | ~P3_PHYADDRPOINTER_REG_29__SCAN_IN | ~P3_PHYADDRPOINTER_REG_27__SCAN_IN | ~P3_PHYADDRPOINTER_REG_26__SCAN_IN | ~new_n3450_ | ~P3_PHYADDRPOINTER_REG_25__SCAN_IN);
  assign new_n3450_ = P3_PHYADDRPOINTER_REG_24__SCAN_IN & P3_PHYADDRPOINTER_REG_22__SCAN_IN & P3_PHYADDRPOINTER_REG_23__SCAN_IN & P3_PHYADDRPOINTER_REG_21__SCAN_IN & new_n3452_ & P3_PHYADDRPOINTER_REG_1__SCAN_IN & new_n3451_ & P3_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign new_n3451_ = P3_PHYADDRPOINTER_REG_15__SCAN_IN & P3_PHYADDRPOINTER_REG_14__SCAN_IN & P3_PHYADDRPOINTER_REG_13__SCAN_IN & P3_PHYADDRPOINTER_REG_12__SCAN_IN & P3_PHYADDRPOINTER_REG_11__SCAN_IN & new_n3302_ & new_n3303_;
  assign new_n3452_ = P3_PHYADDRPOINTER_REG_19__SCAN_IN & P3_PHYADDRPOINTER_REG_20__SCAN_IN & P3_PHYADDRPOINTER_REG_17__SCAN_IN & P3_PHYADDRPOINTER_REG_18__SCAN_IN;
  assign new_n3453_ = new_n3461_ & ((new_n3450_ ^ P3_PHYADDRPOINTER_REG_25__SCAN_IN) ^ (new_n3454_ & ~new_n3459_ & (new_n3450_ | new_n3460_)));
  assign new_n3454_ = ~new_n3458_ & ~new_n3455_ & new_n3456_;
  assign new_n3455_ = (P3_PHYADDRPOINTER_REG_16__SCAN_IN | (new_n3451_ & P3_PHYADDRPOINTER_REG_1__SCAN_IN)) & (~P3_PHYADDRPOINTER_REG_1__SCAN_IN | ~new_n3451_ | ~P3_PHYADDRPOINTER_REG_16__SCAN_IN);
  assign new_n3456_ = (P3_PHYADDRPOINTER_REG_15__SCAN_IN | ~P3_PHYADDRPOINTER_REG_1__SCAN_IN | ~P3_PHYADDRPOINTER_REG_14__SCAN_IN | ~P3_PHYADDRPOINTER_REG_13__SCAN_IN | ~P3_PHYADDRPOINTER_REG_12__SCAN_IN | ~new_n3301_ | ~P3_PHYADDRPOINTER_REG_11__SCAN_IN) & (~P3_PHYADDRPOINTER_REG_15__SCAN_IN | (P3_PHYADDRPOINTER_REG_1__SCAN_IN & P3_PHYADDRPOINTER_REG_14__SCAN_IN & P3_PHYADDRPOINTER_REG_13__SCAN_IN & P3_PHYADDRPOINTER_REG_12__SCAN_IN & new_n3301_ & P3_PHYADDRPOINTER_REG_11__SCAN_IN)) & ((P3_PHYADDRPOINTER_REG_1__SCAN_IN & P3_PHYADDRPOINTER_REG_14__SCAN_IN & P3_PHYADDRPOINTER_REG_13__SCAN_IN & P3_PHYADDRPOINTER_REG_12__SCAN_IN & new_n3301_ & P3_PHYADDRPOINTER_REG_11__SCAN_IN) | (~P3_PHYADDRPOINTER_REG_14__SCAN_IN & (~P3_PHYADDRPOINTER_REG_1__SCAN_IN | ~P3_PHYADDRPOINTER_REG_13__SCAN_IN | ~P3_PHYADDRPOINTER_REG_12__SCAN_IN | ~new_n3301_ | ~P3_PHYADDRPOINTER_REG_11__SCAN_IN))) & (P3_PHYADDRPOINTER_REG_14__SCAN_IN | (~P3_PHYADDRPOINTER_REG_13__SCAN_IN & (~P3_PHYADDRPOINTER_REG_12__SCAN_IN | ~P3_PHYADDRPOINTER_REG_11__SCAN_IN | ~new_n3301_ | ~P3_PHYADDRPOINTER_REG_1__SCAN_IN))) & new_n3457_ & (P3_PHYADDRPOINTER_REG_11__SCAN_IN | ~new_n3301_ | ~P3_PHYADDRPOINTER_REG_1__SCAN_IN) & (~P3_PHYADDRPOINTER_REG_11__SCAN_IN | (new_n3301_ & P3_PHYADDRPOINTER_REG_1__SCAN_IN)) & (~P3_PHYADDRPOINTER_REG_12__SCAN_IN ^ (P3_PHYADDRPOINTER_REG_11__SCAN_IN & new_n3301_ & P3_PHYADDRPOINTER_REG_1__SCAN_IN));
  assign new_n3457_ = P3_PHYADDRPOINTER_REG_10__SCAN_IN & new_n3334_ & P3_PHYADDRPOINTER_REG_9__SCAN_IN & P3_PHYADDRPOINTER_REG_7__SCAN_IN & P3_PHYADDRPOINTER_REG_8__SCAN_IN & ~P3_PHYADDRPOINTER_REG_0__SCAN_IN & P3_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign new_n3458_ = (P3_PHYADDRPOINTER_REG_1__SCAN_IN & new_n3451_ & P3_PHYADDRPOINTER_REG_16__SCAN_IN) ? (~P3_PHYADDRPOINTER_REG_19__SCAN_IN | ~P3_PHYADDRPOINTER_REG_20__SCAN_IN | ~P3_PHYADDRPOINTER_REG_17__SCAN_IN | ~P3_PHYADDRPOINTER_REG_18__SCAN_IN) : (P3_PHYADDRPOINTER_REG_17__SCAN_IN | P3_PHYADDRPOINTER_REG_18__SCAN_IN | P3_PHYADDRPOINTER_REG_19__SCAN_IN | P3_PHYADDRPOINTER_REG_20__SCAN_IN);
  assign new_n3459_ = P3_PHYADDRPOINTER_REG_21__SCAN_IN ^ (new_n3452_ & P3_PHYADDRPOINTER_REG_1__SCAN_IN & new_n3451_ & P3_PHYADDRPOINTER_REG_16__SCAN_IN);
  assign new_n3460_ = ~P3_PHYADDRPOINTER_REG_24__SCAN_IN & ~P3_PHYADDRPOINTER_REG_22__SCAN_IN & ~P3_PHYADDRPOINTER_REG_23__SCAN_IN & (~P3_PHYADDRPOINTER_REG_21__SCAN_IN | ~new_n3452_ | ~P3_PHYADDRPOINTER_REG_1__SCAN_IN | ~new_n3451_ | ~P3_PHYADDRPOINTER_REG_16__SCAN_IN);
  assign new_n3461_ = (((~new_n3334_ | P3_PHYADDRPOINTER_REG_0__SCAN_IN | ~P3_PHYADDRPOINTER_REG_1__SCAN_IN) & (~new_n3334_ | ~P3_PHYADDRPOINTER_REG_7__SCAN_IN) & (new_n3334_ | P3_PHYADDRPOINTER_REG_7__SCAN_IN)) | (new_n3334_ & P3_PHYADDRPOINTER_REG_7__SCAN_IN & ~P3_PHYADDRPOINTER_REG_0__SCAN_IN & P3_PHYADDRPOINTER_REG_1__SCAN_IN)) & P3_PHYADDRPOINTER_REG_3__SCAN_IN & (P3_PHYADDRPOINTER_REG_0__SCAN_IN ^ P3_PHYADDRPOINTER_REG_1__SCAN_IN);
  assign new_n3462_ = P3_PHYADDRPOINTER_REG_26__SCAN_IN & new_n3450_ & P3_PHYADDRPOINTER_REG_25__SCAN_IN;
  assign new_n3463_ = (~P3_PHYADDRPOINTER_REG_26__SCAN_IN ^ (new_n3450_ & P3_PHYADDRPOINTER_REG_25__SCAN_IN)) & (new_n3450_ ^ ~P3_PHYADDRPOINTER_REG_25__SCAN_IN) & (new_n3450_ | new_n3460_) & ~new_n3459_ & ~new_n3458_ & ~new_n3455_ & new_n3456_;
  assign new_n3464_ = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign new_n3465_ = new_n3501_ & new_n3503_ & new_n3466_ & ~new_n3491_ & ~new_n3496_;
  assign new_n3466_ = (~new_n3467_ | new_n3490_) & (new_n3469_ | new_n3470_ | ~new_n3475_ | (~new_n3471_ & P3_EBX_REG_27__SCAN_IN));
  assign new_n3467_ = ~P1_STATE2_REG_0__SCAN_IN & (new_n3312_ | (new_n3468_ & new_n2567_ & (new_n2478_ | new_n2482_)));
  assign new_n3468_ = new_n2495_ & (new_n2585_ | (new_n2529_ & new_n2509_));
  assign new_n3469_ = new_n3449_ & ~new_n3444_ & P3_STATE2_REG_1__SCAN_IN & (~new_n3463_ | (new_n3462_ ^ P3_PHYADDRPOINTER_REG_27__SCAN_IN)) & (new_n3463_ | (new_n3462_ & P3_PHYADDRPOINTER_REG_27__SCAN_IN) | (~new_n3462_ & ~P3_PHYADDRPOINTER_REG_27__SCAN_IN));
  assign new_n3470_ = (~new_n3462_ | ~P3_PHYADDRPOINTER_REG_27__SCAN_IN) & (new_n3462_ | P3_PHYADDRPOINTER_REG_27__SCAN_IN) & ~new_n3449_ & ~new_n3444_ & P3_STATE2_REG_1__SCAN_IN;
  assign new_n3471_ = (P3_EBX_REG_31__SCAN_IN | new_n3474_ | ~new_n3473_ | new_n3444_ | ~P3_STATE2_REG_2__SCAN_IN) & ((new_n3474_ & new_n2947_) | ~new_n3472_ | new_n3444_ | ~P3_STATE2_REG_2__SCAN_IN);
  assign new_n3472_ = new_n2802_ & ~new_n2809_;
  assign new_n3473_ = ~new_n2802_ & ~new_n2809_;
  assign new_n3474_ = ~new_n2943_ & ~P3_STATEBS16_REG_SCAN_IN;
  assign new_n3475_ = (~new_n3476_ | ~new_n3477_) & (new_n3483_ | (new_n3484_ & P3_REIP_REG_27__SCAN_IN) | (~new_n3484_ & ~P3_REIP_REG_27__SCAN_IN)) & (~new_n3444_ | ~P3_REIP_REG_27__SCAN_IN) & (~P3_PHYADDRPOINTER_REG_27__SCAN_IN | new_n3444_ | ~P3_STATE2_REG_3__SCAN_IN);
  assign new_n3476_ = P3_EBX_REG_31__SCAN_IN & ~new_n3474_ & new_n3473_ & P3_STATE2_REG_2__SCAN_IN & (~new_n3448_ | (new_n3445_ & ~new_n3447_));
  assign new_n3477_ = ~P3_EBX_REG_27__SCAN_IN ^ (~P3_EBX_REG_26__SCAN_IN & ~P3_EBX_REG_25__SCAN_IN & new_n3478_ & new_n3482_);
  assign new_n3478_ = ~P3_EBX_REG_21__SCAN_IN & ~P3_EBX_REG_16__SCAN_IN & new_n3479_ & new_n3481_ & ~P3_EBX_REG_17__SCAN_IN & ~P3_EBX_REG_18__SCAN_IN & ~P3_EBX_REG_19__SCAN_IN & ~P3_EBX_REG_20__SCAN_IN;
  assign new_n3479_ = ~P3_EBX_REG_10__SCAN_IN & ~P3_EBX_REG_9__SCAN_IN & new_n3480_ & ~P3_EBX_REG_8__SCAN_IN;
  assign new_n3480_ = ~P3_EBX_REG_7__SCAN_IN & ~P3_EBX_REG_6__SCAN_IN & ~P3_EBX_REG_4__SCAN_IN & ~P3_EBX_REG_5__SCAN_IN & ~P3_EBX_REG_3__SCAN_IN & ~P3_EBX_REG_2__SCAN_IN & ~P3_EBX_REG_0__SCAN_IN & ~P3_EBX_REG_1__SCAN_IN;
  assign new_n3481_ = ~P3_EBX_REG_11__SCAN_IN & ~P3_EBX_REG_12__SCAN_IN & ~P3_EBX_REG_15__SCAN_IN & ~P3_EBX_REG_13__SCAN_IN & ~P3_EBX_REG_14__SCAN_IN;
  assign new_n3482_ = ~P3_EBX_REG_24__SCAN_IN & ~P3_EBX_REG_22__SCAN_IN & ~P3_EBX_REG_23__SCAN_IN;
  assign new_n3483_ = (~new_n3474_ | ~new_n2947_ | ~new_n3472_ | ~P3_STATE2_REG_2__SCAN_IN | (new_n3448_ & (~new_n3445_ | new_n3447_))) & (~new_n3474_ | ~new_n3473_ | ~P3_STATE2_REG_2__SCAN_IN | (new_n3448_ & (~new_n3445_ | new_n3447_)));
  assign new_n3484_ = new_n3485_ & P3_REIP_REG_25__SCAN_IN & P3_REIP_REG_26__SCAN_IN;
  assign new_n3485_ = new_n3489_ & P3_REIP_REG_21__SCAN_IN & new_n3488_ & P3_REIP_REG_16__SCAN_IN & new_n3487_ & P3_REIP_REG_10__SCAN_IN & new_n3486_ & P3_REIP_REG_9__SCAN_IN;
  assign new_n3486_ = P3_REIP_REG_8__SCAN_IN & P3_REIP_REG_7__SCAN_IN & P3_REIP_REG_3__SCAN_IN & P3_REIP_REG_1__SCAN_IN & P3_REIP_REG_2__SCAN_IN & P3_REIP_REG_6__SCAN_IN & P3_REIP_REG_4__SCAN_IN & P3_REIP_REG_5__SCAN_IN;
  assign new_n3487_ = P3_REIP_REG_11__SCAN_IN & P3_REIP_REG_12__SCAN_IN & P3_REIP_REG_15__SCAN_IN & P3_REIP_REG_13__SCAN_IN & P3_REIP_REG_14__SCAN_IN;
  assign new_n3488_ = P3_REIP_REG_19__SCAN_IN & P3_REIP_REG_20__SCAN_IN & P3_REIP_REG_17__SCAN_IN & P3_REIP_REG_18__SCAN_IN;
  assign new_n3489_ = P3_REIP_REG_24__SCAN_IN & P3_REIP_REG_22__SCAN_IN & P3_REIP_REG_23__SCAN_IN;
  assign new_n3490_ = ~P1_UWORD_REG_6__SCAN_IN & ~P1_UWORD_REG_7__SCAN_IN & ~P1_UWORD_REG_2__SCAN_IN & ~P1_UWORD_REG_4__SCAN_IN & ~P1_UWORD_REG_11__SCAN_IN & ~P1_LWORD_REG_7__SCAN_IN & ~P1_LWORD_REG_14__SCAN_IN & ~P1_LWORD_REG_15__SCAN_IN;
  assign new_n3491_ = ((new_n3454_ & ~new_n3459_) | (~new_n3454_ & new_n3459_) | ~new_n3449_ | new_n3444_ | ~P3_STATE2_REG_1__SCAN_IN) & new_n3492_ & (new_n3471_ | ~P3_EBX_REG_21__SCAN_IN) & (~new_n3459_ | new_n3449_ | new_n3444_ | ~P3_STATE2_REG_1__SCAN_IN);
  assign new_n3492_ = (~new_n3476_ | ~new_n3495_) & (~new_n3444_ | ~P3_REIP_REG_21__SCAN_IN) & (~P3_PHYADDRPOINTER_REG_21__SCAN_IN | new_n3444_ | ~P3_STATE2_REG_3__SCAN_IN) & (new_n3483_ | (new_n3493_ & P3_REIP_REG_21__SCAN_IN) | (~new_n3493_ & ~P3_REIP_REG_21__SCAN_IN));
  assign new_n3493_ = new_n3488_ & new_n3494_ & P3_REIP_REG_16__SCAN_IN;
  assign new_n3494_ = new_n3487_ & P3_REIP_REG_10__SCAN_IN & new_n3486_ & P3_REIP_REG_9__SCAN_IN;
  assign new_n3495_ = ~P3_EBX_REG_21__SCAN_IN ^ (~P3_EBX_REG_16__SCAN_IN & new_n3479_ & new_n3481_ & ~P3_EBX_REG_17__SCAN_IN & ~P3_EBX_REG_18__SCAN_IN & ~P3_EBX_REG_19__SCAN_IN & ~P3_EBX_REG_20__SCAN_IN);
  assign new_n3496_ = ((new_n3455_ & ~new_n3456_) | (~new_n3455_ & new_n3456_) | ~new_n3449_ | new_n3444_ | ~P3_STATE2_REG_1__SCAN_IN) & new_n3497_ & (new_n3471_ | ~P3_EBX_REG_16__SCAN_IN) & (~new_n3455_ | new_n3449_ | new_n3444_ | ~P3_STATE2_REG_1__SCAN_IN);
  assign new_n3497_ = (~new_n3476_ | ~new_n3500_) & new_n3499_ & (~new_n3498_ | ~P3_PHYADDRPOINTER_REG_16__SCAN_IN) & (new_n3483_ | (new_n3494_ & P3_REIP_REG_16__SCAN_IN) | (~new_n3494_ & ~P3_REIP_REG_16__SCAN_IN));
  assign new_n3498_ = P3_STATE2_REG_3__SCAN_IN & (~new_n3448_ | (new_n3445_ & ~new_n3447_));
  assign new_n3499_ = (new_n3448_ & (~new_n3445_ | new_n3447_)) ? ~P3_REIP_REG_16__SCAN_IN : (P3_STATE2_REG_1__SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN);
  assign new_n3500_ = ~P3_EBX_REG_16__SCAN_IN ^ (new_n3479_ & new_n3481_);
  assign new_n3501_ = (~new_n3502_ | (~P1_REIP_REG_29__SCAN_IN & ~P1_REIP_REG_12__SCAN_IN)) & ((new_n3425_ & P3_INSTADDRPOINTER_REG_12__SCAN_IN) | ~new_n3307_ | (~new_n3425_ & ~P3_INSTADDRPOINTER_REG_12__SCAN_IN));
  assign new_n3502_ = ~P1_STATE2_REG_2__SCAN_IN & ~P1_STATE2_REG_1__SCAN_IN & (new_n2606_ | (new_n2605_ & ~new_n2073_ & (new_n2478_ | new_n2482_)));
  assign new_n3503_ = (new_n3504_ | new_n3506_) & ((new_n3349_ & new_n2509_) | (~P1_LWORD_REG_11__SCAN_IN & ~P1_LWORD_REG_8__SCAN_IN & ~P1_LWORD_REG_9__SCAN_IN));
  assign new_n3504_ = ~P1_STATE2_REG_0__SCAN_IN & (new_n2997_ | (P1_STATE2_REG_3__SCAN_IN & (new_n2478_ | new_n2482_))) & ~new_n3505_ & (new_n3353_ | ~P1_STATE2_REG_3__SCAN_IN);
  assign new_n3505_ = P1_STATE2_REG_2__SCAN_IN & (~new_n2120_ | ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  assign new_n3506_ = ~P1_INSTQUEUE_REG_14__5__SCAN_IN & ~P1_INSTQUEUE_REG_14__0__SCAN_IN;
  assign new_n3507_ = new_n3512_ & new_n3515_ & new_n3508_ & ~new_n3511_ & (~new_n3086_ | new_n1322_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n3508_ = (new_n3510_ | ~new_n3509_ | ~new_n2114_) & (new_n3509_ | new_n3312_ | (~P1_DATAO_REG_7__SCAN_IN & ~P1_DATAO_REG_15__SCAN_IN & ~P1_DATAO_REG_14__SCAN_IN));
  assign new_n3509_ = new_n3468_ & new_n2567_ & (new_n2478_ | new_n2482_);
  assign new_n3510_ = ~P1_EAX_REG_27__SCAN_IN & ~P1_EAX_REG_23__SCAN_IN & ~P1_EAX_REG_18__SCAN_IN & ~P1_EAX_REG_22__SCAN_IN & ~P1_EAX_REG_20__SCAN_IN;
  assign new_n3511_ = ~new_n3509_ & ~new_n3312_ & (P1_DATAO_REG_27__SCAN_IN | P1_DATAO_REG_23__SCAN_IN | P1_DATAO_REG_18__SCAN_IN | P1_DATAO_REG_22__SCAN_IN | P1_DATAO_REG_20__SCAN_IN);
  assign new_n3512_ = (new_n3513_ | new_n2724_ | ~P2_STATE2_REG_3__SCAN_IN) & (new_n3514_ | new_n2604_ | new_n2606_);
  assign new_n3513_ = ~P2_PHYADDRPOINTER_REG_13__SCAN_IN & ~P2_PHYADDRPOINTER_REG_15__SCAN_IN & ~P2_PHYADDRPOINTER_REG_20__SCAN_IN & ~P2_PHYADDRPOINTER_REG_22__SCAN_IN & ~P2_PHYADDRPOINTER_REG_25__SCAN_IN & ~P2_PHYADDRPOINTER_REG_31__SCAN_IN;
  assign new_n3514_ = ~P1_PHYADDRPOINTER_REG_12__SCAN_IN & ~P1_PHYADDRPOINTER_REG_6__SCAN_IN & ~P1_PHYADDRPOINTER_REG_29__SCAN_IN & ~P1_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign new_n3515_ = (new_n3516_ | new_n3523_) & (new_n3530_ | (new_n2495_ & ((new_n2106_ & new_n2494_) | (new_n2477_ & new_n2493_))));
  assign new_n3516_ = (~P3_STATE2_REG_0__SCAN_IN | ~P3_STATE2_REG_2__SCAN_IN | P3_STATE2_REG_1__SCAN_IN | (~new_n3517_ & new_n3519_ & new_n3521_)) & (P3_STATE2_REG_0__SCAN_IN ? (~P3_FLUSH_REG_SCAN_IN | ~P3_STATE2_REG_2__SCAN_IN | ~P3_STATE2_REG_1__SCAN_IN) : ~P3_STATE2_REG_3__SCAN_IN);
  assign new_n3517_ = new_n2942_ & new_n2947_ & (new_n2840_ | new_n3518_);
  assign new_n3518_ = new_n2802_ & new_n2815_ & ~new_n2826_ & ~new_n2821_ & new_n2796_ & ~new_n2809_ & new_n2790_ & new_n2833_;
  assign new_n3519_ = (new_n3520_ | ~new_n2942_) & (~new_n2853_ | ~new_n2945_);
  assign new_n3520_ = new_n2802_ ? (~new_n2833_ | new_n2790_ | new_n2796_ | new_n2826_ | ~new_n2821_ | ~new_n2809_ | new_n2815_) : (~new_n2815_ | new_n2826_ | new_n2821_ | ~new_n2796_ | new_n2809_ | ~new_n2790_ | ~new_n2833_);
  assign new_n3521_ = new_n2948_ & (~new_n2854_ | ~new_n2945_) & (new_n3522_ | ~new_n2815_ | new_n2833_);
  assign new_n3522_ = new_n2790_ & ~new_n2796_;
  assign new_n3523_ = (new_n3524_ | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_1__SCAN_IN) & (~new_n3529_ | ~P3_STATE2_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) & (~P3_STATE2_REG_1__SCAN_IN | ~P3_INSTADDRPOINTER_REG_0__SCAN_IN | (P3_INSTADDRPOINTER_REG_1__SCAN_IN ^ P3_INSTADDRPOINTER_REG_31__SCAN_IN));
  assign new_n3524_ = (P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | (new_n3527_ & ((~new_n2789_ & new_n3526_) | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN))) & (~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | (~new_n3525_ & new_n3526_)) & (~new_n2832_ | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (new_n3528_ | (P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) | (~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN));
  assign new_n3525_ = new_n2826_ & new_n2833_ & new_n2802_ & new_n2809_ & new_n2815_ & new_n2821_ & ~new_n2790_ & new_n2796_;
  assign new_n3526_ = (~new_n2815_ | ((~new_n2802_ | new_n2809_ | (~new_n2821_ & (~new_n2790_ | new_n2796_) & ~new_n2826_ & (new_n2790_ | ~new_n2796_))) & (~new_n2809_ | ((~new_n2790_ | ~new_n2833_) & (~new_n2802_ | new_n2790_ | new_n2796_))) & ((new_n2796_ & new_n2826_) | new_n2802_ | (~new_n2826_ & ~new_n2821_)))) & (new_n2796_ | ~new_n2821_ | (new_n2809_ & (~new_n2802_ | ~new_n2826_))) & (new_n2796_ | new_n2802_ | ~new_n2790_ | ~new_n2833_) & (new_n2802_ | ~new_n2790_ | ~new_n2826_) & ((~new_n2790_ & ~new_n2796_) | new_n2802_ | ~new_n2809_) & (~new_n2796_ | new_n2821_ | (new_n2790_ & new_n2833_)) & (new_n2833_ | ((~new_n2802_ | new_n2809_) & ~new_n2826_ & (new_n2790_ | new_n2796_))) & (new_n2815_ | (new_n2821_ & (new_n2790_ ? new_n2826_ : ~new_n2796_))) & (~new_n2790_ | ~new_n2821_ | ((~new_n2802_ | ~new_n2809_ | new_n2826_ | ~new_n2815_ | new_n2833_) & (~new_n2826_ | ~new_n2833_ | ~new_n2796_ | new_n2815_))) & (new_n2802_ | new_n2809_ | ~new_n2826_ | ~new_n2833_ | ~new_n2815_ | ~new_n2821_ | new_n2790_ | ~new_n2796_) & (~new_n2826_ | ~new_n2821_ | ~new_n2833_ | new_n2790_ | new_n2796_ | new_n2815_ | new_n2802_ | ~new_n2809_) & (new_n2802_ | ~new_n2833_ | new_n2790_ | new_n2796_ | ~new_n2815_ | new_n2826_ | new_n2821_);
  assign new_n3527_ = (~new_n2815_ | new_n2826_ | new_n2821_ | ~new_n2796_ | new_n2809_ | ~new_n2790_ | ~new_n2833_) & (new_n2826_ | ~new_n2821_ | ~new_n2833_ | new_n2790_ | new_n2796_ | new_n2815_ | new_n2802_ | ~new_n2809_) & (new_n2826_ | ~new_n2802_ | ~new_n2809_ | ~new_n2815_ | ~new_n2821_ | new_n2790_ | ~new_n2796_);
  assign new_n3528_ = (~new_n2790_ | new_n2796_ | ~new_n2802_ | ~new_n2809_ | new_n2826_ | ~new_n2815_ | new_n2833_) & (new_n2802_ | new_n2809_ | new_n2826_ | new_n2821_ | ~new_n2790_ | new_n2796_ | ~new_n2815_ | new_n2833_);
  assign new_n3529_ = P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign new_n3530_ = ~P1_EBX_REG_19__SCAN_IN & ~P1_EBX_REG_23__SCAN_IN & ~P1_EBX_REG_20__SCAN_IN;
  assign new_n3531_ = new_n3532_ & new_n3534_ & new_n3536_ & (~new_n3537_ | new_n1317_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN) & (~new_n3538_ | new_n1317_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n3532_ = (~new_n3370_ | new_n1350_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN) & ((~new_n2666_ & ~new_n3374_) ? P2_READREQUEST_REG_SCAN_IN : ~new_n3533_);
  assign new_n3533_ = P2_STATE2_REG_2__SCAN_IN & (~new_n1322_ ^ ~new_n1370_);
  assign new_n3534_ = (~new_n3201_ | new_n1345_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN) & (new_n3535_ | ~new_n1759_ | ~new_n1330_ | new_n1335_);
  assign new_n3535_ = new_n3078_ & (new_n2976_ | ~BUF2_REG_6__SCAN_IN) & (~new_n2976_ | ~BUF1_REG_6__SCAN_IN) & (new_n2976_ | ~BUF2_REG_14__SCAN_IN) & (~new_n2976_ | ~BUF1_REG_14__SCAN_IN);
  assign new_n3536_ = (~new_n3062_ | new_n1370_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN) & (~new_n3381_ | new_n1345_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n3537_ = new_n3127_ & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n3538_ = ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & new_n3364_ & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n3539_ = new_n3540_ & (new_n3194_ | new_n1317_ | ~new_n1759_ | new_n1335_) & (new_n3544_ | (~new_n1330_ & new_n1317_) | ~new_n1759_ | new_n1335_) & (new_n3090_ | new_n1317_ | ~new_n1759_ | new_n1335_);
  assign new_n3540_ = (new_n1759_ | new_n3541_) & (~new_n2724_ | new_n3542_) & (~new_n3439_ | ~new_n3543_) & (~new_n2724_ | (~P2_REIP_REG_13__SCAN_IN & ~P2_REIP_REG_15__SCAN_IN));
  assign new_n3541_ = ~P2_EAX_REG_10__SCAN_IN & ~P2_EAX_REG_13__SCAN_IN & ~P2_EAX_REG_14__SCAN_IN & ~P2_EAX_REG_21__SCAN_IN & ~P2_EAX_REG_22__SCAN_IN & ~P2_EAX_REG_30__SCAN_IN;
  assign new_n3542_ = ~P2_REIP_REG_25__SCAN_IN & ~P2_REIP_REG_31__SCAN_IN & ~P2_REIP_REG_20__SCAN_IN & ~P2_REIP_REG_22__SCAN_IN;
  assign new_n3543_ = P2_STATE2_REG_0__SCAN_IN & (P2_EAX_REG_7__SCAN_IN | P2_EAX_REG_10__SCAN_IN);
  assign new_n3544_ = (~new_n2976_ | ~BUF1_REG_14__SCAN_IN) & (new_n2976_ | ~BUF2_REG_14__SCAN_IN) & (~new_n2976_ | ~BUF1_REG_10__SCAN_IN) & (new_n2976_ | ~BUF2_REG_10__SCAN_IN) & (~new_n2976_ | ~BUF1_REG_13__SCAN_IN) & (new_n2976_ | ~BUF2_REG_13__SCAN_IN);
  assign new_n3545_ = new_n3986_ & new_n3546_ & new_n3924_ & new_n3936_ & new_n3907_ & new_n3556_ & new_n3578_;
  assign new_n3546_ = ~new_n3547_ & (~P2_FLUSH_REG_SCAN_IN | (~new_n3554_ & new_n1791_)) & (new_n2683_ | (~P2_EBX_REG_31__SCAN_IN & ~P2_EBX_REG_5__SCAN_IN & ~P2_EBX_REG_24__SCAN_IN));
  assign new_n3547_ = (~P3_REIP_REG_2__SCAN_IN | P3_STATE2_REG_2__SCAN_IN | (~new_n2937_ & ~new_n3282_)) & (~P3_INSTADDRPOINTER_REG_2__SCAN_IN | new_n2937_ | new_n3282_) & (~new_n2937_ | (~new_n3548_ & ~new_n3549_ & new_n3550_));
  assign new_n3548_ = (new_n2850_ | (~new_n2844_ & ~new_n2849_)) & (~new_n2857_ | ~new_n2860_ | new_n2859_ | new_n2846_ | new_n2844_ | new_n2849_);
  assign new_n3549_ = ((new_n2883_ & ~P3_INSTADDRPOINTER_REG_0__SCAN_IN & (new_n2873_ | ~P3_INSTADDRPOINTER_REG_1__SCAN_IN)) | (~new_n2873_ & ~new_n2883_) | (new_n2873_ & ~P3_INSTADDRPOINTER_REG_1__SCAN_IN) | (~P3_INSTADDRPOINTER_REG_2__SCAN_IN & (new_n2867_ | new_n2873_ | new_n2883_) & (~new_n2867_ | (~new_n2873_ & ~new_n2883_))) | (P3_INSTADDRPOINTER_REG_2__SCAN_IN & (new_n2867_ ^ (~new_n2873_ & ~new_n2883_)))) & new_n2928_ & (((~new_n2883_ | P3_INSTADDRPOINTER_REG_0__SCAN_IN | (~new_n2873_ & P3_INSTADDRPOINTER_REG_1__SCAN_IN)) & (new_n2873_ | new_n2883_) & (~new_n2873_ | P3_INSTADDRPOINTER_REG_1__SCAN_IN)) | (~P3_INSTADDRPOINTER_REG_2__SCAN_IN ^ (~new_n2867_ ^ (~new_n2873_ & ~new_n2883_))));
  assign new_n3550_ = ((new_n3552_ & (new_n3551_ | P3_INSTADDRPOINTER_REG_2__SCAN_IN) & (~new_n3551_ | ~P3_INSTADDRPOINTER_REG_2__SCAN_IN)) | ~new_n2927_ | (~new_n3552_ & (new_n3551_ ^ ~P3_INSTADDRPOINTER_REG_2__SCAN_IN))) & (~new_n2858_ | (P3_INSTADDRPOINTER_REG_2__SCAN_IN & P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN) | (~P3_INSTADDRPOINTER_REG_2__SCAN_IN & (~P3_INSTADDRPOINTER_REG_0__SCAN_IN | ~P3_INSTADDRPOINTER_REG_1__SCAN_IN))) & (new_n3553_ | (P3_INSTADDRPOINTER_REG_1__SCAN_IN & P3_INSTADDRPOINTER_REG_2__SCAN_IN) | (~P3_INSTADDRPOINTER_REG_1__SCAN_IN & ~P3_INSTADDRPOINTER_REG_2__SCAN_IN));
  assign new_n3551_ = new_n2867_ ^ new_n2873_;
  assign new_n3552_ = (new_n2873_ | P3_INSTADDRPOINTER_REG_1__SCAN_IN) & (new_n2919_ | (new_n2873_ & P3_INSTADDRPOINTER_REG_1__SCAN_IN));
  assign new_n3553_ = (new_n2826_ | ~new_n2802_ | ~new_n2809_ | ~new_n2815_ | ~new_n2821_ | new_n2790_ | ~new_n2796_) & (~new_n2833_ | new_n2790_ | new_n2796_ | new_n2826_ | ~new_n2821_ | ~new_n2809_ | new_n2815_) & (~new_n2815_ | new_n2826_ | new_n2821_ | ~new_n2796_ | new_n2809_ | ~new_n2790_ | ~new_n2833_);
  assign new_n3554_ = new_n3555_ & (new_n1322_ | ~new_n1370_ | (~new_n1762_ & (new_n1768_ | ~new_n1781_)));
  assign new_n3555_ = (new_n1788_ | (~new_n1322_ & new_n1370_)) & (new_n1786_ | (new_n1787_ & ~new_n1370_)) & (new_n1790_ | (~new_n2670_ & (~new_n1322_ | ~new_n1370_) & (new_n1322_ | new_n1370_)));
  assign new_n3556_ = new_n3562_ & new_n3564_ & new_n3557_ & new_n3560_ & new_n3566_ & (~new_n3516_ | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n3557_ = (new_n3293_ | ~new_n3297_ | (~new_n3455_ & ~new_n3558_)) & (new_n3559_ | new_n3293_ | ~new_n3284_);
  assign new_n3558_ = P3_PHYADDRPOINTER_REG_12__SCAN_IN ^ (P3_PHYADDRPOINTER_REG_11__SCAN_IN & new_n3301_ & P3_PHYADDRPOINTER_REG_1__SCAN_IN);
  assign new_n3559_ = ~P3_REIP_REG_16__SCAN_IN & ~P3_REIP_REG_21__SCAN_IN & ~P3_REIP_REG_0__SCAN_IN & ~P3_REIP_REG_12__SCAN_IN;
  assign new_n3560_ = (~new_n3561_ | ((~P3_PHYADDRPOINTER_REG_21__SCAN_IN | (new_n3452_ & new_n3451_ & P3_PHYADDRPOINTER_REG_16__SCAN_IN)) & (~new_n3300_ ^ P3_PHYADDRPOINTER_REG_12__SCAN_IN) & (P3_PHYADDRPOINTER_REG_21__SCAN_IN | ~new_n3452_ | ~new_n3451_ | ~P3_PHYADDRPOINTER_REG_16__SCAN_IN))) & (~new_n3561_ | (~P3_PHYADDRPOINTER_REG_0__SCAN_IN & (~new_n3451_ ^ P3_PHYADDRPOINTER_REG_16__SCAN_IN)));
  assign new_n3561_ = new_n3305_ & (new_n3294_ | (new_n2950_ & ((new_n2927_ & new_n2939_) | (new_n2928_ & new_n2945_))));
  assign new_n3562_ = (~new_n3498_ | new_n3563_) & (~P3_PHYADDRPOINTER_REG_0__SCAN_IN | new_n3293_ | ~new_n3297_);
  assign new_n3563_ = ~P3_PHYADDRPOINTER_REG_1__SCAN_IN & ~P3_PHYADDRPOINTER_REG_3__SCAN_IN & ~P3_PHYADDRPOINTER_REG_7__SCAN_IN & ~P3_PHYADDRPOINTER_REG_10__SCAN_IN & ~P3_PHYADDRPOINTER_REG_25__SCAN_IN & ~P3_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign new_n3564_ = (~new_n3558_ | new_n3293_ | ~new_n3298_) & (new_n3565_ | (~P3_EAX_REG_21__SCAN_IN & ~P3_EAX_REG_5__SCAN_IN & ~P3_EAX_REG_8__SCAN_IN));
  assign new_n3565_ = new_n2950_ & (new_n3525_ | (new_n2853_ & new_n2945_) | (~new_n3520_ & new_n2942_));
  assign new_n3566_ = new_n3567_ & ~new_n3576_ & ((~new_n3455_ & ~P3_PHYADDRPOINTER_REG_0__SCAN_IN) | new_n3293_ | ~new_n3298_);
  assign new_n3567_ = (new_n2950_ & (new_n3525_ | (~new_n3520_ & new_n2942_) | (new_n2853_ & new_n2945_))) ? ~new_n3568_ : new_n3575_;
  assign new_n3568_ = new_n2826_ & ((~P3_EAX_REG_28__SCAN_IN & new_n3574_ & P3_EAX_REG_23__SCAN_IN & P3_EAX_REG_22__SCAN_IN & new_n3569_ & P3_EAX_REG_21__SCAN_IN) | (P3_EAX_REG_28__SCAN_IN & (~new_n3574_ | ~P3_EAX_REG_23__SCAN_IN | ~P3_EAX_REG_22__SCAN_IN | ~new_n3569_ | ~P3_EAX_REG_21__SCAN_IN)) | (P3_EAX_REG_23__SCAN_IN ^ (P3_EAX_REG_22__SCAN_IN & new_n3569_ & P3_EAX_REG_21__SCAN_IN)) | ~new_n3573_ | (new_n3569_ ^ P3_EAX_REG_21__SCAN_IN));
  assign new_n3569_ = new_n3571_ & new_n3572_ & P3_EAX_REG_9__SCAN_IN & P3_EAX_REG_10__SCAN_IN & new_n3570_ & P3_EAX_REG_8__SCAN_IN;
  assign new_n3570_ = P3_EAX_REG_6__SCAN_IN & P3_EAX_REG_7__SCAN_IN & P3_EAX_REG_5__SCAN_IN & P3_EAX_REG_0__SCAN_IN & P3_EAX_REG_1__SCAN_IN & P3_EAX_REG_4__SCAN_IN & P3_EAX_REG_2__SCAN_IN & P3_EAX_REG_3__SCAN_IN;
  assign new_n3571_ = P3_EAX_REG_19__SCAN_IN & P3_EAX_REG_20__SCAN_IN & P3_EAX_REG_17__SCAN_IN & P3_EAX_REG_18__SCAN_IN;
  assign new_n3572_ = P3_EAX_REG_11__SCAN_IN & P3_EAX_REG_12__SCAN_IN & P3_EAX_REG_13__SCAN_IN & P3_EAX_REG_14__SCAN_IN & P3_EAX_REG_15__SCAN_IN & P3_EAX_REG_16__SCAN_IN;
  assign new_n3573_ = (~new_n3570_ ^ P3_EAX_REG_8__SCAN_IN) & (~P3_EAX_REG_5__SCAN_IN ^ (P3_EAX_REG_0__SCAN_IN & P3_EAX_REG_1__SCAN_IN & P3_EAX_REG_4__SCAN_IN & P3_EAX_REG_2__SCAN_IN & P3_EAX_REG_3__SCAN_IN));
  assign new_n3574_ = P3_EAX_REG_26__SCAN_IN & P3_EAX_REG_27__SCAN_IN & P3_EAX_REG_24__SCAN_IN & P3_EAX_REG_25__SCAN_IN;
  assign new_n3575_ = ~P3_EAX_REG_23__SCAN_IN & ~P3_EAX_REG_28__SCAN_IN;
  assign new_n3576_ = new_n3577_ & P3_STATE2_REG_2__SCAN_IN & (~new_n3448_ | (new_n3445_ & ~new_n3447_));
  assign new_n3577_ = new_n2809_ & ((P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN & (~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN)) | (~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) | (~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN));
  assign new_n3578_ = new_n3888_ & new_n3902_ & new_n3830_ & new_n3822_ & new_n3580_ & ~new_n3579_ & new_n3587_ & new_n3784_;
  assign new_n3579_ = ~new_n3444_ & ~P3_STATE2_REG_1__SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN;
  assign new_n3580_ = new_n3584_ & (~new_n3583_ | ~P3_EAX_REG_10__SCAN_IN) & (~P3_MORE_REG_SCAN_IN | (~new_n3581_ & new_n2950_));
  assign new_n3581_ = ~new_n3582_ & new_n3446_ & (new_n2943_ | (~new_n2947_ & (~new_n2802_ ^ new_n2815_)));
  assign new_n3582_ = (~new_n2796_ | new_n2809_ | ~new_n2790_ | ~new_n2833_ | ~new_n2815_ | new_n2826_ | new_n2821_) & (~new_n2833_ | new_n2790_ | new_n2796_ | new_n2826_ | ~new_n2821_ | ~new_n2809_ | new_n2815_);
  assign new_n3583_ = new_n3445_ & new_n2947_ & (new_n2840_ | new_n3518_);
  assign new_n3584_ = (new_n3585_ | ~P2_LWORD_REG_15__SCAN_IN) & (~new_n3440_ | ~P2_EAX_REG_15__SCAN_IN);
  assign new_n3585_ = new_n1340_ & ~new_n3586_ & new_n1792_ & new_n1788_ & new_n1350_ & new_n1356_ & new_n1330_ & new_n1377_;
  assign new_n3586_ = new_n1790_ & (~new_n1325_ | ~new_n1326_ | ~new_n1323_ | ~new_n1324_);
  assign new_n3587_ = ~new_n3755_ & new_n3757_ & new_n3728_ & new_n3749_ & new_n3588_ & new_n3608_;
  assign new_n3588_ = new_n3603_ & ~new_n3594_ & ((new_n3596_ & ~new_n2821_ & new_n3602_) | ~new_n3589_ | (~new_n3595_ & P3_INSTQUEUE_REG_0__3__SCAN_IN));
  assign new_n3589_ = new_n3590_ & (~new_n3592_ | ~BUF2_REG_3__SCAN_IN | new_n3593_ | (P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) | (~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)));
  assign new_n3590_ = (~new_n3591_ | ~BUF2_REG_27__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (~new_n3591_ | ~BUF2_REG_19__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  assign new_n3591_ = P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (~P3_STATE2_REG_2__SCAN_IN ^ ~P3_STATE2_REG_1__SCAN_IN));
  assign new_n3592_ = ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (~P3_STATE2_REG_2__SCAN_IN ^ ~P3_STATE2_REG_1__SCAN_IN));
  assign new_n3593_ = (~P3_STATEBS16_REG_SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN) & ~P3_STATE2_REG_2__SCAN_IN & (P3_STATEBS16_REG_SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN);
  assign new_n3594_ = new_n3598_ & (new_n3595_ | ~P3_INSTQUEUE_REG_0__4__SCAN_IN) & (~new_n3596_ | new_n2833_ | ~new_n3602_);
  assign new_n3595_ = ~new_n3597_ & new_n3592_ & (new_n3596_ | ~P3_STATE2_REG_3__SCAN_IN);
  assign new_n3596_ = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3597_ = ((~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))) & (P3_STATE2_REG_2__SCAN_IN | (~P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN) | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN));
  assign new_n3598_ = (~new_n3599_ | new_n3593_ | (P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) | (~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))) & (~new_n3600_ | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (~new_n3601_ | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  assign new_n3599_ = BUF2_REG_4__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (P3_STATE2_REG_2__SCAN_IN ^ P3_STATE2_REG_1__SCAN_IN));
  assign new_n3600_ = BUF2_REG_28__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (P3_STATE2_REG_2__SCAN_IN ^ P3_STATE2_REG_1__SCAN_IN)) & P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN;
  assign new_n3601_ = BUF2_REG_20__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (P3_STATE2_REG_2__SCAN_IN ^ P3_STATE2_REG_1__SCAN_IN)) & P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN;
  assign new_n3602_ = P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (~P3_STATE2_REG_2__SCAN_IN ^ ~P3_STATE2_REG_1__SCAN_IN));
  assign new_n3603_ = ((P2_DATAO_REG_20__SCAN_IN & ~new_n3604_ & new_n3606_) | (new_n3604_ & P1_DATAO_REG_20__SCAN_IN) | (BUF1_REG_20__SCAN_IN & ~new_n3604_ & ~new_n3606_)) & ((P2_DATAO_REG_7__SCAN_IN & ~new_n3604_ & new_n3606_) | (new_n3604_ & P1_DATAO_REG_7__SCAN_IN) | (BUF1_REG_7__SCAN_IN & ~new_n3604_ & ~new_n3606_));
  assign new_n3604_ = new_n3605_ & P1_ADDRESS_REG_29__SCAN_IN & (~new_n2957_ | ~new_n2958_ | ~new_n2955_ | ~new_n2956_);
  assign new_n3605_ = ~P1_BE_N_REG_3__SCAN_IN & ~P1_BE_N_REG_2__SCAN_IN & ~P1_BE_N_REG_1__SCAN_IN & ~P1_BE_N_REG_0__SCAN_IN & ~P1_ADS_N_REG_SCAN_IN & P1_M_IO_N_REG_SCAN_IN & ~P1_D_C_N_REG_SCAN_IN & P1_W_R_N_REG_SCAN_IN;
  assign new_n3606_ = new_n3607_ & P2_ADDRESS_REG_29__SCAN_IN & (~new_n2979_ | ~new_n2980_ | ~new_n2977_ | ~new_n2978_);
  assign new_n3607_ = ~P2_BE_N_REG_1__SCAN_IN & ~P2_BE_N_REG_0__SCAN_IN & ~P2_BE_N_REG_3__SCAN_IN & ~P2_BE_N_REG_2__SCAN_IN & P2_W_R_N_REG_SCAN_IN & ~P2_D_C_N_REG_SCAN_IN & P2_M_IO_N_REG_SCAN_IN & ~P2_ADS_N_REG_SCAN_IN;
  assign new_n3608_ = new_n3711_ & new_n3717_ & new_n3726_ & new_n3609_ & new_n3687_ & new_n3634_ & new_n3670_ & new_n3679_;
  assign new_n3609_ = new_n3615_ & new_n3610_ & new_n3611_ & new_n3626_ & new_n3619_ & new_n3623_;
  assign new_n3610_ = (~new_n3591_ | ~BUF2_REG_19__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (~new_n3591_ | ~BUF2_REG_23__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  assign new_n3611_ = (~new_n3612_ | ~new_n3614_) & (~P3_STATE_REG_2__SCAN_IN | (new_n3613_ & ((P3_STATE_REG_0__SCAN_IN ? (P3_STATE_REG_2__SCAN_IN | ~P3_STATE_REG_1__SCAN_IN) : P3_STATE_REG_1__SCAN_IN) ? P3_STATEBS16_REG_SCAN_IN : BS16)));
  assign new_n3612_ = BUF2_REG_27__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (P3_STATE2_REG_2__SCAN_IN ^ P3_STATE2_REG_1__SCAN_IN)) & P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN;
  assign new_n3613_ = (~P3_STATE_REG_1__SCAN_IN | (~HOLD & (~READY2 | ~READY22_REG_SCAN_IN))) & (~HOLD | ~P3_STATE_REG_0__SCAN_IN) & (NA | P3_STATE_REG_0__SCAN_IN);
  assign new_n3614_ = P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3615_ = (~new_n3601_ | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (~new_n3616_ | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (~new_n3617_ | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (~new_n3618_ | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  assign new_n3616_ = BUF2_REG_31__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (P3_STATE2_REG_2__SCAN_IN ^ P3_STATE2_REG_1__SCAN_IN)) & P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN;
  assign new_n3617_ = BUF2_REG_24__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (P3_STATE2_REG_2__SCAN_IN ^ P3_STATE2_REG_1__SCAN_IN)) & P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN;
  assign new_n3618_ = BUF2_REG_22__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (P3_STATE2_REG_2__SCAN_IN ^ P3_STATE2_REG_1__SCAN_IN)) & P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN;
  assign new_n3619_ = (~new_n3620_ | ~new_n3622_) & (~P3_INSTQUEUE_REG_9__1__SCAN_IN | (new_n3592_ & ~new_n3621_));
  assign new_n3620_ = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3621_ = ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_STATEBS16_REG_SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN);
  assign new_n3622_ = BUF2_REG_29__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (P3_STATE2_REG_2__SCAN_IN ^ P3_STATE2_REG_1__SCAN_IN)) & P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN;
  assign new_n3623_ = (~new_n3625_ | ~new_n3591_ | ~BUF2_REG_19__SCAN_IN) & (~new_n3624_ | ~new_n3591_ | ~BUF2_REG_31__SCAN_IN);
  assign new_n3624_ = P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3625_ = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3626_ = (~new_n3630_ | ~new_n3631_) & (~new_n3599_ | ~new_n3629_) & (~new_n3632_ | ~new_n3633_) & (~new_n3628_ | (~new_n3627_ & ~new_n3632_));
  assign new_n3627_ = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n3628_ = BUF2_REG_23__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (P3_STATE2_REG_2__SCAN_IN ^ P3_STATE2_REG_1__SCAN_IN)) & P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN;
  assign new_n3629_ = ((P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN) | P3_STATE2_REG_2__SCAN_IN | (~P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN)) & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN));
  assign new_n3630_ = P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n3631_ = BUF2_REG_16__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (P3_STATE2_REG_2__SCAN_IN ^ P3_STATE2_REG_1__SCAN_IN)) & P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN;
  assign new_n3632_ = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3633_ = BUF2_REG_30__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (P3_STATE2_REG_2__SCAN_IN ^ P3_STATE2_REG_1__SCAN_IN)) & P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN;
  assign new_n3634_ = new_n3642_ & new_n3635_ & new_n3639_ & new_n3661_ & new_n3656_ & new_n3659_ & new_n3648_ & new_n3651_;
  assign new_n3635_ = ~new_n3637_ & (~new_n3636_ | (P3_ADDRESS_REG_15__SCAN_IN & P3_ADDRESS_REG_20__SCAN_IN & ~P3_ADDRESS_REG_16__SCAN_IN)) & ~new_n3638_ & (new_n3636_ | (P2_ADDRESS_REG_28__SCAN_IN & P2_ADDRESS_REG_17__SCAN_IN));
  assign new_n3636_ = (P1_DATAO_REG_31__SCAN_IN | ~P1_DATAO_REG_30__SCAN_IN) & (~P2_DATAO_REG_30__SCAN_IN | P2_DATAO_REG_31__SCAN_IN) & (~P3_DATAO_REG_30__SCAN_IN | P3_DATAO_REG_31__SCAN_IN);
  assign new_n3637_ = P2_STATE2_REG_1__SCAN_IN & ((~P2_STATE2_REG_0__SCAN_IN & P2_STATEBS16_REG_SCAN_IN) | ((~READY12_REG_SCAN_IN | ~READY21_REG_SCAN_IN) & ~P2_STATE2_REG_2__SCAN_IN & P2_STATE2_REG_0__SCAN_IN));
  assign new_n3638_ = (P1_DATAWIDTH_REG_30__SCAN_IN | P1_DATAWIDTH_REG_24__SCAN_IN | P1_DATAWIDTH_REG_26__SCAN_IN) & (P1_STATE_REG_1__SCAN_IN | P1_STATE_REG_0__SCAN_IN) & (~P1_STATE_REG_0__SCAN_IN | P1_STATE_REG_2__SCAN_IN | ~P1_STATE_REG_1__SCAN_IN);
  assign new_n3639_ = ~new_n3640_ & ~new_n3641_ & (~new_n3636_ | (P3_ADDRESS_REG_28__SCAN_IN & P3_ADDRESS_REG_17__SCAN_IN)) & (new_n3636_ | (~P2_ADDRESS_REG_21__SCAN_IN & ~P2_ADDRESS_REG_16__SCAN_IN));
  assign new_n3640_ = (HOLD | P3_REQUESTPENDING_REG_SCAN_IN) & (P3_STATE_REG_1__SCAN_IN | ~P3_REQUESTPENDING_REG_SCAN_IN) & ~P3_STATE_REG_2__SCAN_IN & P3_STATE_REG_0__SCAN_IN & (~P3_STATE_REG_1__SCAN_IN | (READY2 & READY22_REG_SCAN_IN)) & (~NA | P3_STATE_REG_2__SCAN_IN | ~P3_STATE_REG_1__SCAN_IN);
  assign new_n3641_ = (P1_DATAWIDTH_REG_5__SCAN_IN | P1_DATAWIDTH_REG_9__SCAN_IN) & (P1_STATE_REG_1__SCAN_IN | P1_STATE_REG_0__SCAN_IN) & (~P1_STATE_REG_0__SCAN_IN | P1_STATE_REG_2__SCAN_IN | ~P1_STATE_REG_1__SCAN_IN);
  assign new_n3642_ = ~new_n3644_ & ~new_n3645_ & ~new_n3646_ & ~new_n3647_ & (~new_n3643_ | ~new_n3592_ | ~BUF2_REG_5__SCAN_IN);
  assign new_n3643_ = P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ((P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN) | P3_STATE2_REG_2__SCAN_IN | (~P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN));
  assign new_n3644_ = (~P1_STATE_REG_1__SCAN_IN | P1_STATE_REG_0__SCAN_IN) & (P1_BE_N_REG_1__SCAN_IN | P1_ADDRESS_REG_29__SCAN_IN | P1_ADDRESS_REG_7__SCAN_IN | P1_ADDRESS_REG_24__SCAN_IN | P1_ADDRESS_REG_9__SCAN_IN);
  assign new_n3645_ = (P1_STATE_REG_2__SCAN_IN | ~P1_REIP_REG_29__SCAN_IN | ~P1_REIP_REG_17__SCAN_IN) & P1_STATE_REG_1__SCAN_IN & ~P1_STATE_REG_0__SCAN_IN & (~P1_STATE_REG_2__SCAN_IN | ~P1_REIP_REG_28__SCAN_IN | ~P1_REIP_REG_16__SCAN_IN);
  assign new_n3646_ = (P1_STATE_REG_2__SCAN_IN | ~P1_REIP_REG_12__SCAN_IN | P1_REIP_REG_11__SCAN_IN) & P1_STATE_REG_1__SCAN_IN & ~P1_STATE_REG_0__SCAN_IN & (~P1_STATE_REG_2__SCAN_IN | ~P1_REIP_REG_11__SCAN_IN | P1_REIP_REG_8__SCAN_IN);
  assign new_n3647_ = ~P3_STATE_REG_2__SCAN_IN & P3_STATE_REG_1__SCAN_IN & ~P3_STATE_REG_0__SCAN_IN & (P3_REIP_REG_4__SCAN_IN | P3_REIP_REG_14__SCAN_IN | P3_REIP_REG_29__SCAN_IN | P3_REIP_REG_17__SCAN_IN | P3_REIP_REG_22__SCAN_IN);
  assign new_n3648_ = new_n3650_ & new_n3649_ & (P1_STATE_REG_1__SCAN_IN | P1_STATE_REG_0__SCAN_IN) & (~P1_STATE_REG_0__SCAN_IN | P1_STATE_REG_2__SCAN_IN | ~P1_STATE_REG_1__SCAN_IN);
  assign new_n3649_ = P3_DATAWIDTH_REG_19__SCAN_IN & P3_DATAWIDTH_REG_22__SCAN_IN & P3_DATAWIDTH_REG_23__SCAN_IN & P3_DATAWIDTH_REG_26__SCAN_IN & P3_DATAWIDTH_REG_7__SCAN_IN & P3_DATAWIDTH_REG_9__SCAN_IN & (~P2_STATE2_REG_2__SCAN_IN | P2_STATE2_REG_1__SCAN_IN);
  assign new_n3650_ = (P3_STATE_REG_1__SCAN_IN | P3_STATE_REG_0__SCAN_IN) & (~P3_STATE_REG_0__SCAN_IN | P3_STATE_REG_2__SCAN_IN | ~P3_STATE_REG_1__SCAN_IN) & (P2_STATE_REG_1__SCAN_IN | P2_STATE_REG_0__SCAN_IN) & (~P2_STATE_REG_0__SCAN_IN | P2_STATE_REG_2__SCAN_IN | ~P2_STATE_REG_1__SCAN_IN);
  assign new_n3651_ = new_n3654_ & new_n3655_ & new_n3652_ & new_n3653_;
  assign new_n3652_ = ((P1_STATE_REG_1__SCAN_IN & ~P1_STATE_REG_0__SCAN_IN) | (P1_M_IO_N_REG_SCAN_IN & ~P1_BE_N_REG_0__SCAN_IN)) & ((P2_STATE_REG_1__SCAN_IN & ~P2_STATE_REG_0__SCAN_IN) | (P2_BE_N_REG_3__SCAN_IN & ~P2_ADDRESS_REG_26__SCAN_IN));
  assign new_n3653_ = (P1_STATE_REG_2__SCAN_IN | P1_STATE_REG_1__SCAN_IN | P1_STATE_REG_0__SCAN_IN) & ((~P2_STATE_REG_2__SCAN_IN & P2_BYTEENABLE_REG_3__SCAN_IN) | ~P2_STATE_REG_1__SCAN_IN | P2_STATE_REG_0__SCAN_IN);
  assign new_n3654_ = P2_DATAWIDTH_REG_13__SCAN_IN & P2_DATAWIDTH_REG_17__SCAN_IN & P3_DATAWIDTH_REG_28__SCAN_IN & P2_DATAWIDTH_REG_7__SCAN_IN & P1_DATAWIDTH_REG_12__SCAN_IN & P2_DATAWIDTH_REG_23__SCAN_IN & P2_DATAWIDTH_REG_28__SCAN_IN;
  assign new_n3655_ = (~P3_MEMORYFETCH_REG_SCAN_IN | ~P3_STATE_REG_1__SCAN_IN | P3_STATE_REG_0__SCAN_IN) & (~P2_CODEFETCH_REG_SCAN_IN | ~P2_STATE_REG_1__SCAN_IN | P2_STATE_REG_0__SCAN_IN);
  assign new_n3656_ = new_n3657_ & ~new_n3658_ & (~P2_REIP_REG_27__SCAN_IN | ~P2_STATE_REG_2__SCAN_IN | ~P2_STATE_REG_1__SCAN_IN | P2_STATE_REG_0__SCAN_IN);
  assign new_n3657_ = ((~P3_REIP_REG_3__SCAN_IN & ~P3_REIP_REG_5__SCAN_IN) | P3_STATE_REG_2__SCAN_IN | ~P3_STATE_REG_1__SCAN_IN | P3_STATE_REG_0__SCAN_IN) & ((P3_STATE_REG_1__SCAN_IN & ~P3_STATE_REG_0__SCAN_IN) | (~P3_ADDRESS_REG_15__SCAN_IN & ~P3_ADDRESS_REG_27__SCAN_IN & ~P3_ADDRESS_REG_20__SCAN_IN));
  assign new_n3658_ = P1_STATE_REG_2__SCAN_IN & P1_STATE_REG_1__SCAN_IN & ~P1_STATE_REG_0__SCAN_IN & (P1_REIP_REG_10__SCAN_IN | P1_REIP_REG_30__SCAN_IN | P1_REIP_REG_25__SCAN_IN);
  assign new_n3659_ = new_n3660_ & (~P1_STATE_REG_1__SCAN_IN | P1_STATE_REG_0__SCAN_IN | (~P1_BYTEENABLE_REG_1__SCAN_IN & P1_MEMORYFETCH_REG_SCAN_IN & ~P1_BYTEENABLE_REG_0__SCAN_IN)) & (~P1_REIP_REG_9__SCAN_IN | P1_STATE_REG_2__SCAN_IN | ~P1_STATE_REG_1__SCAN_IN | P1_STATE_REG_0__SCAN_IN);
  assign new_n3660_ = (~P3_REIP_REG_2__SCAN_IN | ~P3_STATE_REG_2__SCAN_IN | ~P3_STATE_REG_1__SCAN_IN | P3_STATE_REG_0__SCAN_IN) & (P2_D_C_N_REG_SCAN_IN | (~P2_STATE_REG_0__SCAN_IN & (~P2_STATE_REG_2__SCAN_IN | P2_STATE_REG_1__SCAN_IN)));
  assign new_n3661_ = new_n3664_ & ~new_n3662_ & ~new_n3663_ & ~new_n3668_ & ~new_n3669_ & ~new_n3665_ & ~new_n3666_ & new_n3667_;
  assign new_n3662_ = (P3_STATE_REG_1__SCAN_IN & ~P3_STATE_REG_0__SCAN_IN) ? P3_STATE_REG_2__SCAN_IN : (P3_ADDRESS_REG_1__SCAN_IN | P3_ADDRESS_REG_3__SCAN_IN | P3_ADDRESS_REG_2__SCAN_IN);
  assign new_n3663_ = ~P2_ADDRESS_REG_29__SCAN_IN & ((~P1_DATAO_REG_31__SCAN_IN & P1_DATAO_REG_30__SCAN_IN) | (P2_DATAO_REG_30__SCAN_IN & ~P2_DATAO_REG_31__SCAN_IN) | (P3_DATAO_REG_30__SCAN_IN & ~P3_DATAO_REG_31__SCAN_IN));
  assign new_n3664_ = (P3_ADDRESS_REG_29__SCAN_IN | (~P1_DATAO_REG_31__SCAN_IN & P1_DATAO_REG_30__SCAN_IN) | (P3_DATAO_REG_30__SCAN_IN & ~P3_DATAO_REG_31__SCAN_IN) | (P2_DATAO_REG_30__SCAN_IN & ~P2_DATAO_REG_31__SCAN_IN)) & (~P3_ADDRESS_REG_21__SCAN_IN | (~P1_DATAO_REG_31__SCAN_IN & P1_DATAO_REG_30__SCAN_IN) | (P3_DATAO_REG_30__SCAN_IN & ~P3_DATAO_REG_31__SCAN_IN) | (P2_DATAO_REG_30__SCAN_IN & ~P2_DATAO_REG_31__SCAN_IN));
  assign new_n3665_ = (P1_DATAWIDTH_REG_16__SCAN_IN | P1_DATAWIDTH_REG_1__SCAN_IN | P1_DATAWIDTH_REG_14__SCAN_IN) & (P1_STATE_REG_1__SCAN_IN | P1_STATE_REG_0__SCAN_IN) & (~P1_STATE_REG_0__SCAN_IN | P1_STATE_REG_2__SCAN_IN | ~P1_STATE_REG_1__SCAN_IN);
  assign new_n3666_ = ~P1_ADDRESS_REG_10__SCAN_IN & (~P1_STATE_REG_1__SCAN_IN | P1_STATE_REG_0__SCAN_IN);
  assign new_n3667_ = ((P3_STATE_REG_1__SCAN_IN & ~P3_STATE_REG_0__SCAN_IN) | (~P3_ADDRESS_REG_12__SCAN_IN & ~P3_M_IO_N_REG_SCAN_IN)) & ((P1_STATE_REG_1__SCAN_IN & ~P1_STATE_REG_0__SCAN_IN) | (P1_ADDRESS_REG_27__SCAN_IN & P1_ADDRESS_REG_15__SCAN_IN));
  assign new_n3668_ = (P3_DATAWIDTH_REG_31__SCAN_IN | P3_DATAWIDTH_REG_10__SCAN_IN | P3_DATAWIDTH_REG_17__SCAN_IN) & (P3_STATE_REG_1__SCAN_IN | P3_STATE_REG_0__SCAN_IN) & (~P3_STATE_REG_0__SCAN_IN | P3_STATE_REG_2__SCAN_IN | ~P3_STATE_REG_1__SCAN_IN);
  assign new_n3669_ = (~P2_ADDRESS_REG_20__SCAN_IN | ~P2_ADDRESS_REG_15__SCAN_IN) & ((~P1_DATAO_REG_31__SCAN_IN & P1_DATAO_REG_30__SCAN_IN) | (P2_DATAO_REG_30__SCAN_IN & ~P2_DATAO_REG_31__SCAN_IN) | (P3_DATAO_REG_30__SCAN_IN & ~P3_DATAO_REG_31__SCAN_IN));
  assign new_n3670_ = ~new_n3671_ & (new_n3672_ | P3_BYTEENABLE_REG_3__SCAN_IN) & ~new_n3677_ & (~new_n3672_ | (~P3_DATAWIDTH_REG_1__SCAN_IN & (~P3_REIP_REG_1__SCAN_IN | (~P3_DATAWIDTH_REG_0__SCAN_IN & ~P3_REIP_REG_0__SCAN_IN))));
  assign new_n3671_ = new_n3591_ & BUF2_REG_17__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n3672_ = new_n3675_ & new_n3676_ & new_n3673_ & new_n3674_;
  assign new_n3673_ = ~P3_DATAWIDTH_REG_18__SCAN_IN & ~P3_DATAWIDTH_REG_19__SCAN_IN & ~P3_DATAWIDTH_REG_15__SCAN_IN & ~P3_DATAWIDTH_REG_16__SCAN_IN & ~P3_DATAWIDTH_REG_20__SCAN_IN & ~P3_DATAWIDTH_REG_21__SCAN_IN & ~P3_DATAWIDTH_REG_22__SCAN_IN & ~P3_DATAWIDTH_REG_23__SCAN_IN;
  assign new_n3674_ = ~P3_DATAWIDTH_REG_26__SCAN_IN & ~P3_DATAWIDTH_REG_27__SCAN_IN & ~P3_DATAWIDTH_REG_24__SCAN_IN & ~P3_DATAWIDTH_REG_25__SCAN_IN & ~P3_DATAWIDTH_REG_28__SCAN_IN & ~P3_DATAWIDTH_REG_29__SCAN_IN & ~P3_DATAWIDTH_REG_30__SCAN_IN & ~P3_DATAWIDTH_REG_31__SCAN_IN;
  assign new_n3675_ = ~P3_DATAWIDTH_REG_2__SCAN_IN & ~P3_DATAWIDTH_REG_3__SCAN_IN & ~P3_DATAWIDTH_REG_4__SCAN_IN & ~P3_DATAWIDTH_REG_5__SCAN_IN & (~P3_DATAWIDTH_REG_0__SCAN_IN | ~P3_DATAWIDTH_REG_1__SCAN_IN) & ~P3_DATAWIDTH_REG_10__SCAN_IN & ~P3_DATAWIDTH_REG_17__SCAN_IN;
  assign new_n3676_ = ~P3_DATAWIDTH_REG_8__SCAN_IN & ~P3_DATAWIDTH_REG_9__SCAN_IN & ~P3_DATAWIDTH_REG_6__SCAN_IN & ~P3_DATAWIDTH_REG_7__SCAN_IN & ~P3_DATAWIDTH_REG_11__SCAN_IN & ~P3_DATAWIDTH_REG_12__SCAN_IN & ~P3_DATAWIDTH_REG_13__SCAN_IN & ~P3_DATAWIDTH_REG_14__SCAN_IN;
  assign new_n3677_ = (new_n3607_ & ~P2_ADDRESS_REG_29__SCAN_IN) ? ~new_n3678_ : (BUF2_REG_18__SCAN_IN | ~BUF2_REG_1__SCAN_IN | BUF2_REG_10__SCAN_IN);
  assign new_n3678_ = ~P2_DATAO_REG_6__SCAN_IN & ~P2_DATAO_REG_10__SCAN_IN & ~P2_DATAO_REG_14__SCAN_IN & P2_DATAO_REG_24__SCAN_IN;
  assign new_n3679_ = new_n3685_ & (new_n3680_ | ~P2_BYTEENABLE_REG_3__SCAN_IN) & ((~P3_STATE_REG_1__SCAN_IN & ~P3_STATE_REG_0__SCAN_IN) | (BS16 & (P3_STATE_REG_0__SCAN_IN ? (~P3_STATE_REG_2__SCAN_IN & P3_STATE_REG_1__SCAN_IN) : ~P3_STATE_REG_1__SCAN_IN)) | (P3_STATEBS16_REG_SCAN_IN & (P3_STATE_REG_1__SCAN_IN | P3_STATE_REG_0__SCAN_IN) & (~P3_STATE_REG_0__SCAN_IN | P3_STATE_REG_2__SCAN_IN | ~P3_STATE_REG_1__SCAN_IN)));
  assign new_n3680_ = new_n3683_ & new_n3684_ & new_n3681_ & new_n3682_;
  assign new_n3681_ = ~P2_DATAWIDTH_REG_18__SCAN_IN & ~P2_DATAWIDTH_REG_19__SCAN_IN & ~P2_DATAWIDTH_REG_16__SCAN_IN & ~P2_DATAWIDTH_REG_17__SCAN_IN & ~P2_DATAWIDTH_REG_20__SCAN_IN & ~P2_DATAWIDTH_REG_21__SCAN_IN & ~P2_DATAWIDTH_REG_22__SCAN_IN & ~P2_DATAWIDTH_REG_23__SCAN_IN;
  assign new_n3682_ = ~P2_DATAWIDTH_REG_26__SCAN_IN & ~P2_DATAWIDTH_REG_27__SCAN_IN & ~P2_DATAWIDTH_REG_24__SCAN_IN & ~P2_DATAWIDTH_REG_25__SCAN_IN & ~P2_DATAWIDTH_REG_28__SCAN_IN & ~P2_DATAWIDTH_REG_29__SCAN_IN & ~P2_DATAWIDTH_REG_30__SCAN_IN & ~P2_DATAWIDTH_REG_31__SCAN_IN;
  assign new_n3683_ = ~P2_DATAWIDTH_REG_4__SCAN_IN & ~P2_DATAWIDTH_REG_5__SCAN_IN & ~P2_DATAWIDTH_REG_6__SCAN_IN & ~P2_DATAWIDTH_REG_7__SCAN_IN & ~P2_DATAWIDTH_REG_2__SCAN_IN & ~P2_DATAWIDTH_REG_3__SCAN_IN & (~P2_DATAWIDTH_REG_0__SCAN_IN | ~P2_DATAWIDTH_REG_1__SCAN_IN);
  assign new_n3684_ = ~P2_DATAWIDTH_REG_10__SCAN_IN & ~P2_DATAWIDTH_REG_11__SCAN_IN & ~P2_DATAWIDTH_REG_8__SCAN_IN & ~P2_DATAWIDTH_REG_9__SCAN_IN & ~P2_DATAWIDTH_REG_12__SCAN_IN & ~P2_DATAWIDTH_REG_13__SCAN_IN & ~P2_DATAWIDTH_REG_14__SCAN_IN & ~P2_DATAWIDTH_REG_15__SCAN_IN;
  assign new_n3685_ = (~new_n3686_ | ~new_n3592_ | ~BUF2_REG_1__SCAN_IN) & ((P1_STATEBS16_REG_SCAN_IN & (P1_STATE_REG_1__SCAN_IN | P1_STATE_REG_0__SCAN_IN) & (~P1_STATE_REG_0__SCAN_IN | P1_STATE_REG_2__SCAN_IN | ~P1_STATE_REG_1__SCAN_IN)) | (~P1_STATE_REG_2__SCAN_IN & ~P1_STATE_REG_1__SCAN_IN & ~P1_STATE_REG_0__SCAN_IN) | (BS16 & (P1_STATE_REG_0__SCAN_IN ? (~P1_STATE_REG_2__SCAN_IN & P1_STATE_REG_1__SCAN_IN) : ~P1_STATE_REG_1__SCAN_IN)));
  assign new_n3686_ = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ((P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN) | P3_STATE2_REG_2__SCAN_IN | (~P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN));
  assign new_n3687_ = new_n3688_ & new_n3690_ & new_n3704_ & new_n3693_ & new_n3697_ & new_n3702_;
  assign new_n3688_ = (~new_n3643_ | ((~new_n3592_ | ~BUF2_REG_2__SCAN_IN) & (~new_n3592_ | ~BUF2_REG_4__SCAN_IN))) & (~new_n3689_ | ((~new_n3592_ | ~BUF2_REG_1__SCAN_IN) & (~new_n3592_ | ~BUF2_REG_7__SCAN_IN)));
  assign new_n3689_ = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & (P3_STATE2_REG_2__SCAN_IN | (~P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN) | (P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)));
  assign new_n3690_ = (~new_n3600_ | ~new_n3692_) & ((new_n3683_ & new_n3684_ & new_n3681_ & new_n3682_) ? new_n3691_ : P2_BYTEENABLE_REG_2__SCAN_IN);
  assign new_n3691_ = P2_REIP_REG_1__SCAN_IN ? P2_REIP_REG_0__SCAN_IN : (~P2_DATAWIDTH_REG_1__SCAN_IN & (~P2_DATAWIDTH_REG_0__SCAN_IN | ~P2_REIP_REG_0__SCAN_IN));
  assign new_n3692_ = P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3693_ = ~new_n3694_ & ~new_n3695_ & ((new_n3607_ & ~P2_ADDRESS_REG_29__SCAN_IN) | (~BUF2_REG_11__SCAN_IN & ~BUF2_REG_3__SCAN_IN & ~BUF2_REG_14__SCAN_IN)) & (new_n3696_ | ~new_n3607_ | P2_ADDRESS_REG_29__SCAN_IN);
  assign new_n3694_ = (~P2_REIP_REG_5__SCAN_IN | ~P2_STATE_REG_2__SCAN_IN | ~P2_STATE_REG_1__SCAN_IN | P2_STATE_REG_0__SCAN_IN) & (~P2_REIP_REG_6__SCAN_IN | P2_STATE_REG_2__SCAN_IN | ~P2_STATE_REG_1__SCAN_IN | P2_STATE_REG_0__SCAN_IN) & (~P2_ADDRESS_REG_4__SCAN_IN | (P2_STATE_REG_1__SCAN_IN & ~P2_STATE_REG_0__SCAN_IN));
  assign new_n3695_ = (~P3_REIP_REG_10__SCAN_IN | ~P3_STATE_REG_2__SCAN_IN | ~P3_STATE_REG_1__SCAN_IN | P3_STATE_REG_0__SCAN_IN) & (~P3_REIP_REG_11__SCAN_IN | P3_STATE_REG_2__SCAN_IN | ~P3_STATE_REG_1__SCAN_IN | P3_STATE_REG_0__SCAN_IN) & (~P3_ADDRESS_REG_9__SCAN_IN | (P3_STATE_REG_1__SCAN_IN & ~P3_STATE_REG_0__SCAN_IN));
  assign new_n3696_ = ~P2_DATAO_REG_3__SCAN_IN & ~P2_DATAO_REG_11__SCAN_IN & ~P2_DATAO_REG_31__SCAN_IN & ~P2_DATAO_REG_17__SCAN_IN & ~P2_DATAO_REG_18__SCAN_IN;
  assign new_n3697_ = ~new_n3698_ & ~new_n3700_ & ~new_n3701_ & ~new_n3699_ & (~P2_REIP_REG_28__SCAN_IN | P2_STATE_REG_2__SCAN_IN | ~P2_STATE_REG_1__SCAN_IN | P2_STATE_REG_0__SCAN_IN);
  assign new_n3698_ = (P2_STATE_REG_0__SCAN_IN ? (P2_STATE_REG_2__SCAN_IN | ~P2_STATE_REG_1__SCAN_IN) : P2_STATE_REG_1__SCAN_IN) ? (P2_DATAWIDTH_REG_18__SCAN_IN | P2_DATAWIDTH_REG_1__SCAN_IN | P2_DATAWIDTH_REG_6__SCAN_IN) : (BS16 | (~P2_STATE_REG_2__SCAN_IN & ~P2_STATE_REG_1__SCAN_IN));
  assign new_n3699_ = (P1_REIP_REG_31__SCAN_IN | P1_REIP_REG_26__SCAN_IN) & ~P1_STATE_REG_2__SCAN_IN & P1_STATE_REG_1__SCAN_IN & ~P1_STATE_REG_0__SCAN_IN;
  assign new_n3700_ = P3_STATE_REG_2__SCAN_IN & P3_STATE_REG_1__SCAN_IN & ~P3_STATE_REG_0__SCAN_IN & (P3_REIP_REG_28__SCAN_IN | P3_REIP_REG_3__SCAN_IN | P3_REIP_REG_21__SCAN_IN);
  assign new_n3701_ = P3_STATE_REG_2__SCAN_IN & P3_STATE_REG_1__SCAN_IN & ~P3_STATE_REG_0__SCAN_IN & (P3_REIP_REG_16__SCAN_IN | P3_REIP_REG_4__SCAN_IN | P3_REIP_REG_13__SCAN_IN);
  assign new_n3702_ = (new_n3607_ & ~P2_ADDRESS_REG_29__SCAN_IN) ? (P2_DATAO_REG_27__SCAN_IN & P2_DATAO_REG_1__SCAN_IN & P2_DATAO_REG_15__SCAN_IN) : new_n3703_;
  assign new_n3703_ = ~BUF2_REG_6__SCAN_IN & BUF2_REG_15__SCAN_IN & BUF2_REG_27__SCAN_IN & ~BUF2_REG_31__SCAN_IN & ~BUF2_REG_17__SCAN_IN & BUF2_REG_24__SCAN_IN;
  assign new_n3704_ = (~new_n3705_ | new_n3706_) & ~new_n3707_ & ~new_n3708_ & ~new_n3709_ & ~new_n3710_;
  assign new_n3705_ = P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ((P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN) | P3_STATE2_REG_2__SCAN_IN | (~P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN));
  assign new_n3706_ = (~BUF2_REG_5__SCAN_IN | P3_STATE2_REG_0__SCAN_IN | ((~P3_STATE2_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) & (P3_STATE2_REG_2__SCAN_IN ^ ~P3_STATE2_REG_1__SCAN_IN))) & (~BUF2_REG_0__SCAN_IN | P3_STATE2_REG_0__SCAN_IN | ((~P3_STATE2_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) & (P3_STATE2_REG_2__SCAN_IN ^ ~P3_STATE2_REG_1__SCAN_IN)));
  assign new_n3707_ = (~P3_REIP_REG_13__SCAN_IN | P3_STATE_REG_2__SCAN_IN | ~P3_STATE_REG_1__SCAN_IN | P3_STATE_REG_0__SCAN_IN) & (~P3_REIP_REG_12__SCAN_IN | ~P3_STATE_REG_2__SCAN_IN | ~P3_STATE_REG_1__SCAN_IN | P3_STATE_REG_0__SCAN_IN) & (~P3_ADDRESS_REG_11__SCAN_IN | (P3_STATE_REG_1__SCAN_IN & ~P3_STATE_REG_0__SCAN_IN));
  assign new_n3708_ = (~P1_REIP_REG_30__SCAN_IN | P1_STATE_REG_2__SCAN_IN | ~P1_STATE_REG_1__SCAN_IN | P1_STATE_REG_0__SCAN_IN) & (~P1_REIP_REG_29__SCAN_IN | ~P1_STATE_REG_2__SCAN_IN | ~P1_STATE_REG_1__SCAN_IN | P1_STATE_REG_0__SCAN_IN) & (~P1_ADDRESS_REG_28__SCAN_IN | (P1_STATE_REG_1__SCAN_IN & ~P1_STATE_REG_0__SCAN_IN));
  assign new_n3709_ = (~P2_REIP_REG_12__SCAN_IN | P2_STATE_REG_2__SCAN_IN | ~P2_STATE_REG_1__SCAN_IN | P2_STATE_REG_0__SCAN_IN) & (~P2_REIP_REG_11__SCAN_IN | ~P2_STATE_REG_2__SCAN_IN | ~P2_STATE_REG_1__SCAN_IN | P2_STATE_REG_0__SCAN_IN) & (~P2_ADDRESS_REG_10__SCAN_IN | (P2_STATE_REG_1__SCAN_IN & ~P2_STATE_REG_0__SCAN_IN));
  assign new_n3710_ = (~P3_REIP_REG_8__SCAN_IN | P3_STATE_REG_2__SCAN_IN | ~P3_STATE_REG_1__SCAN_IN | P3_STATE_REG_0__SCAN_IN) & (~P3_REIP_REG_7__SCAN_IN | ~P3_STATE_REG_2__SCAN_IN | ~P3_STATE_REG_1__SCAN_IN | P3_STATE_REG_0__SCAN_IN) & (~P3_ADDRESS_REG_6__SCAN_IN | (P3_STATE_REG_1__SCAN_IN & ~P3_STATE_REG_0__SCAN_IN));
  assign new_n3711_ = new_n3712_ & (new_n3715_ | ~new_n3592_ | ~BUF2_REG_7__SCAN_IN) & (new_n3716_ | new_n3604_ | new_n3606_);
  assign new_n3712_ = (~new_n3625_ | (~new_n3622_ & ~new_n3612_ & ~new_n3600_)) & (~new_n3624_ | (new_n3713_ & new_n3714_));
  assign new_n3713_ = (~BUF2_REG_20__SCAN_IN | P3_STATE2_REG_0__SCAN_IN | ((~P3_STATE2_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) & (P3_STATE2_REG_2__SCAN_IN ^ ~P3_STATE2_REG_1__SCAN_IN)) | ~P3_STATEBS16_REG_SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN) & (~BUF2_REG_21__SCAN_IN | P3_STATE2_REG_0__SCAN_IN | ((~P3_STATE2_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) & (P3_STATE2_REG_2__SCAN_IN ^ ~P3_STATE2_REG_1__SCAN_IN)) | ~P3_STATEBS16_REG_SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN);
  assign new_n3714_ = (~BUF2_REG_16__SCAN_IN | P3_STATE2_REG_0__SCAN_IN | ((~P3_STATE2_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) & (P3_STATE2_REG_2__SCAN_IN ^ ~P3_STATE2_REG_1__SCAN_IN)) | ~P3_STATEBS16_REG_SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN) & (~BUF2_REG_18__SCAN_IN | P3_STATE2_REG_0__SCAN_IN | ((~P3_STATE2_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) & (P3_STATE2_REG_2__SCAN_IN ^ ~P3_STATE2_REG_1__SCAN_IN)) | ~P3_STATEBS16_REG_SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN);
  assign new_n3715_ = ((~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) | ((~P3_STATEBS16_REG_SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN) & ~P3_STATE2_REG_2__SCAN_IN & (P3_STATEBS16_REG_SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN))) & (P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (~P3_STATE2_REG_2__SCAN_IN & (P3_STATEBS16_REG_SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN) & (~P3_STATEBS16_REG_SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN | (~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) | (P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN))));
  assign new_n3716_ = ~BUF1_REG_1__SCAN_IN & ~BUF1_REG_2__SCAN_IN & ~BUF1_REG_12__SCAN_IN & ~BUF1_REG_13__SCAN_IN & ~BUF1_REG_23__SCAN_IN & ~BUF1_REG_31__SCAN_IN;
  assign new_n3717_ = new_n3722_ & ~new_n3723_ & ~new_n3724_ & (new_n3718_ | ~P3_INSTQUEUE_REG_9__7__SCAN_IN) & ~new_n3721_ & (new_n3719_ | ~P3_INSTQUEUE_REG_1__1__SCAN_IN);
  assign new_n3718_ = new_n3592_ & ~new_n3621_;
  assign new_n3719_ = ((~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) | (new_n3720_ & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)) & new_n3592_ & (~P3_STATE2_REG_3__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN));
  assign new_n3720_ = ~P3_STATE2_REG_2__SCAN_IN & (P3_STATEBS16_REG_SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN);
  assign new_n3721_ = new_n3643_ & ((new_n3592_ & BUF2_REG_0__SCAN_IN) | (new_n3592_ & BUF2_REG_3__SCAN_IN));
  assign new_n3722_ = (~new_n3591_ | ~BUF2_REG_25__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (~new_n3591_ | ~BUF2_REG_21__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  assign new_n3723_ = ((new_n3592_ & BUF2_REG_2__SCAN_IN) | (new_n3592_ & BUF2_REG_7__SCAN_IN)) & ~new_n3593_ & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  assign new_n3724_ = (~new_n3720_ | (new_n3725_ & (~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN))) & new_n3592_ & BUF2_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  assign new_n3725_ = P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN;
  assign new_n3726_ = (new_n2802_ | ~new_n3602_ | ~new_n3692_) & (new_n3727_ | new_n3604_ | ~new_n3606_);
  assign new_n3727_ = ~P2_DATAO_REG_1__SCAN_IN & ~P2_DATAO_REG_2__SCAN_IN & ~P2_DATAO_REG_12__SCAN_IN & ~P2_DATAO_REG_13__SCAN_IN & ~P2_DATAO_REG_23__SCAN_IN & ~P2_DATAO_REG_31__SCAN_IN;
  assign new_n3728_ = ~new_n3729_ & ~new_n3735_ & ~new_n3741_ & (~new_n3745_ | (new_n3748_ & ~new_n2790_ & new_n3602_));
  assign new_n3729_ = (~new_n3620_ | new_n2790_ | ~new_n3592_ | ~P3_STATE2_REG_3__SCAN_IN) & ~new_n3731_ & new_n3732_ & (~P3_INSTQUEUE_REG_8__6__SCAN_IN | (~new_n3730_ & new_n3592_ & (new_n3620_ | ~P3_STATE2_REG_3__SCAN_IN)));
  assign new_n3730_ = (~new_n3720_ | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & ((P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ^ (~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)));
  assign new_n3731_ = (~new_n3720_ | (new_n3725_ & (P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)))) & new_n3592_ & BUF2_REG_6__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ^ (~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN));
  assign new_n3732_ = (~new_n3618_ | ~new_n3734_) & (~new_n3733_ | ~new_n3633_);
  assign new_n3733_ = P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3734_ = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3735_ = (~new_n3739_ | new_n2815_ | ~new_n3602_) & (~new_n3738_ | ~new_n3740_) & new_n3737_ & (new_n3736_ | ~P3_INSTQUEUE_REG_10__2__SCAN_IN);
  assign new_n3736_ = ((P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) | (new_n3720_ & ((~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)))) & new_n3592_ & (~P3_STATE2_REG_3__SCAN_IN | (~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN));
  assign new_n3737_ = (~new_n3627_ | ~new_n3591_ | ~BUF2_REG_26__SCAN_IN) & (~new_n3620_ | ~new_n3591_ | ~BUF2_REG_18__SCAN_IN);
  assign new_n3738_ = BUF2_REG_2__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (P3_STATE2_REG_2__SCAN_IN ^ P3_STATE2_REG_1__SCAN_IN));
  assign new_n3739_ = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3740_ = P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P3_STATE2_REG_2__SCAN_IN | (~P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN) | (P3_STATEBS16_REG_SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN & (P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)));
  assign new_n3741_ = (~new_n3625_ | new_n2790_ | ~new_n3592_ | ~P3_STATE2_REG_3__SCAN_IN) & ~new_n3743_ & new_n3744_ & (~P3_INSTQUEUE_REG_12__6__SCAN_IN | (~new_n3742_ & new_n3592_ & (new_n3625_ | ~P3_STATE2_REG_3__SCAN_IN)));
  assign new_n3742_ = (~new_n3720_ | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & (~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)));
  assign new_n3743_ = (~new_n3720_ | (new_n3725_ & (~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)))) & new_n3592_ & BUF2_REG_6__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN));
  assign new_n3744_ = (~new_n3618_ | ~new_n3739_) & (~new_n3630_ | ~new_n3633_);
  assign new_n3745_ = (new_n3746_ | ~P3_INSTQUEUE_REG_2__6__SCAN_IN) & new_n3747_ & (~new_n3596_ | ~new_n3618_);
  assign new_n3746_ = ((~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) | (new_n3720_ & (P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ? (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) : (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)))) & new_n3592_ & (~P3_STATE2_REG_3__SCAN_IN | (~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN));
  assign new_n3747_ = (~new_n3633_ | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (~new_n3592_ | ~BUF2_REG_6__SCAN_IN | new_n3593_ | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN));
  assign new_n3748_ = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3749_ = new_n3750_ & ~new_n3751_ & ((new_n3632_ & ~new_n2796_ & new_n3602_) | ~new_n3754_ | (~new_n3753_ & P3_INSTQUEUE_REG_4__5__SCAN_IN));
  assign new_n3750_ = ((P2_DATAO_REG_21__SCAN_IN & ~new_n3604_ & new_n3606_) | (new_n3604_ & P1_DATAO_REG_21__SCAN_IN) | (BUF1_REG_21__SCAN_IN & ~new_n3604_ & ~new_n3606_)) & ((P2_DATAO_REG_19__SCAN_IN & ~new_n3604_ & new_n3606_) | (new_n3604_ & P1_DATAO_REG_19__SCAN_IN) | (BUF1_REG_19__SCAN_IN & ~new_n3604_ & ~new_n3606_));
  assign new_n3751_ = (~new_n3739_ | new_n2833_ | ~new_n3602_) & (new_n3736_ | ~P3_INSTQUEUE_REG_10__4__SCAN_IN) & new_n3752_ & (~new_n3599_ | ~new_n3740_);
  assign new_n3752_ = (~new_n3601_ | ~new_n3620_) & (~new_n3627_ | ~new_n3600_);
  assign new_n3753_ = ((~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))) | (new_n3720_ & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))) & new_n3592_ & (~P3_STATE2_REG_3__SCAN_IN | (~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN));
  assign new_n3754_ = (~new_n3629_ | ~new_n3592_ | ~BUF2_REG_5__SCAN_IN) & (~new_n3692_ | ~BUF2_REG_29__SCAN_IN | ~new_n3592_ | ~new_n3725_) & (~new_n3748_ | ~BUF2_REG_21__SCAN_IN | ~new_n3592_ | ~new_n3725_);
  assign new_n3755_ = new_n3445_ & new_n3518_ & (~new_n3756_ | P3_EAX_REG_29__SCAN_IN | P3_EAX_REG_22__SCAN_IN | P3_EAX_REG_25__SCAN_IN);
  assign new_n3756_ = ~P3_EAX_REG_6__SCAN_IN & ~P3_EAX_REG_9__SCAN_IN & ~P3_EAX_REG_1__SCAN_IN & ~P3_EAX_REG_3__SCAN_IN & ~P3_EAX_REG_10__SCAN_IN & ~P3_EAX_REG_13__SCAN_IN & ~P3_EAX_REG_14__SCAN_IN & ~P3_EAX_REG_18__SCAN_IN;
  assign new_n3757_ = (new_n3758_ | ~new_n3602_) & new_n3759_ & new_n3765_ & new_n3770_ & new_n3775_ & new_n3779_;
  assign new_n3758_ = ((new_n2802_ & new_n2826_) | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (new_n2833_ | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (new_n2821_ | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  assign new_n3759_ = ~new_n3762_ & ~new_n3763_ & ~new_n3760_ & ~new_n3761_;
  assign new_n3760_ = new_n3627_ & new_n3602_ & (~new_n2791_ | ~new_n2792_ | ~new_n2793_ | ~new_n2794_ | ~new_n2795_);
  assign new_n3761_ = (new_n3596_ | new_n3734_) & new_n3602_ & (~new_n2827_ | ~new_n2828_ | ~new_n2829_ | ~new_n2830_ | ~new_n2831_);
  assign new_n3762_ = new_n3614_ & new_n3602_ & (~new_n2810_ | ~new_n2811_ | ~new_n2812_ | ~new_n2813_ | ~new_n2814_);
  assign new_n3763_ = new_n3764_ & new_n3602_ & (~new_n2797_ | ~new_n2798_ | ~new_n2799_ | ~new_n2800_ | ~new_n2801_);
  assign new_n3764_ = P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n3765_ = ~new_n3766_ & (~new_n3604_ | new_n3769_) & (new_n3753_ | ~P3_INSTQUEUE_REG_4__4__SCAN_IN) & (new_n3746_ | (~P3_INSTQUEUE_REG_2__7__SCAN_IN & ~P3_INSTQUEUE_REG_2__2__SCAN_IN));
  assign new_n3766_ = (new_n3768_ | (~new_n3592_ & (new_n3767_ | ~new_n3295_ | ~P3_STATE2_REG_0__SCAN_IN))) & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ((~P3_STATE2_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (new_n3592_ | (~new_n3767_ & new_n3295_ & P3_STATE2_REG_0__SCAN_IN))));
  assign new_n3767_ = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN & ~P3_FLUSH_REG_SCAN_IN & ((~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3768_ = (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ((P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_1__SCAN_IN) & (P3_STATEBS16_REG_SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN))) & (~P3_STATE2_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_STATEBS16_REG_SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN);
  assign new_n3769_ = ~P1_DATAO_REG_31__SCAN_IN & ~P1_DATAO_REG_23__SCAN_IN & ~P1_DATAO_REG_13__SCAN_IN & ~P1_DATAO_REG_12__SCAN_IN & ~P1_DATAO_REG_2__SCAN_IN & ~P1_DATAO_REG_1__SCAN_IN;
  assign new_n3770_ = new_n3773_ & (new_n3604_ | ~new_n3606_) & new_n3771_ & (~new_n3680_ | ~new_n3774_);
  assign new_n3771_ = ~new_n3772_ & (~new_n3592_ | ~BUF2_REG_6__SCAN_IN | new_n3593_ | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  assign new_n3772_ = P2_REQUESTPENDING_REG_SCAN_IN & ((P2_STATE_REG_0__SCAN_IN & ~P2_STATE_REG_2__SCAN_IN & ~P2_STATE_REG_1__SCAN_IN) | (~HOLD & ((P2_STATE_REG_2__SCAN_IN & (~NA | P2_STATE_REG_0__SCAN_IN)) | (P2_STATE_REG_0__SCAN_IN & (~READY12_REG_SCAN_IN | ~READY21_REG_SCAN_IN)))));
  assign new_n3773_ = (~P3_INSTQUEUE_REG_0__7__SCAN_IN | (~new_n3597_ & new_n3592_ & (new_n3596_ | ~P3_STATE2_REG_3__SCAN_IN))) & (~new_n3596_ | ((~BUF2_REG_18__SCAN_IN | ~new_n3592_ | ~new_n3725_) & (~BUF2_REG_23__SCAN_IN | ~new_n3592_ | ~new_n3725_)));
  assign new_n3774_ = ~P2_DATAWIDTH_REG_1__SCAN_IN & (~P2_REIP_REG_1__SCAN_IN | (~P2_DATAWIDTH_REG_0__SCAN_IN & ~P2_REIP_REG_0__SCAN_IN));
  assign new_n3775_ = new_n3777_ & (~P3_INSTQUEUE_REG_7__6__SCAN_IN | (new_n3776_ & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)) & (new_n3778_ | (new_n3776_ & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN));
  assign new_n3776_ = (new_n3720_ | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & new_n3592_ & (~P3_STATE2_REG_3__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN));
  assign new_n3777_ = (~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ((~new_n3591_ | ~BUF2_REG_26__SCAN_IN) & (~new_n3591_ | ~BUF2_REG_31__SCAN_IN))) & (P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ((~new_n3591_ | ~BUF2_REG_25__SCAN_IN) & (~new_n3591_ | ~BUF2_REG_31__SCAN_IN)));
  assign new_n3778_ = ~P3_INSTQUEUE_REG_15__5__SCAN_IN & ~P3_INSTQUEUE_REG_15__4__SCAN_IN & ~P3_INSTQUEUE_REG_15__0__SCAN_IN & ~P3_INSTQUEUE_REG_15__3__SCAN_IN & ~P3_INSTQUEUE_REG_15__2__SCAN_IN;
  assign new_n3779_ = ~new_n3780_ & ~new_n3781_ & ~new_n3782_ & (new_n3783_ | (~P3_INSTQUEUE_REG_11__5__SCAN_IN & ~P3_INSTQUEUE_REG_11__0__SCAN_IN));
  assign new_n3780_ = new_n3625_ & ((new_n3591_ & BUF2_REG_24__SCAN_IN) | (new_n3591_ & BUF2_REG_26__SCAN_IN));
  assign new_n3781_ = P3_INSTQUEUE_REG_6__7__SCAN_IN & (((P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & (~new_n3720_ | (P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ? (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) : (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)))) | ~new_n3592_ | (P3_STATE2_REG_3__SCAN_IN & (P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)));
  assign new_n3782_ = P3_INSTQUEUE_REG_14__3__SCAN_IN & (((~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & (~new_n3720_ | ((~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)))) | ~new_n3592_ | (P3_STATE2_REG_3__SCAN_IN & (P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)));
  assign new_n3783_ = P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & (new_n3720_ | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & new_n3592_ & (~P3_STATE2_REG_3__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN));
  assign new_n3784_ = ~new_n3785_ & new_n3806_ & new_n3810_ & new_n3787_ & new_n3800_;
  assign new_n3785_ = ~new_n3786_ & new_n3445_ & ~new_n2943_ & new_n2839_ & ~new_n2802_;
  assign new_n3786_ = ~BUF2_REG_6__SCAN_IN & ~BUF2_REG_9__SCAN_IN & ~BUF2_REG_10__SCAN_IN & ~BUF2_REG_13__SCAN_IN & ~BUF2_REG_1__SCAN_IN & ~BUF2_REG_2__SCAN_IN & ~BUF2_REG_3__SCAN_IN & ~BUF2_REG_14__SCAN_IN;
  assign new_n3787_ = ~new_n3788_ & ~new_n3790_ & ~new_n3792_ & (~new_n3796_ | (new_n3733_ & ~new_n2809_ & new_n3602_));
  assign new_n3788_ = (~new_n3630_ | new_n2796_ | ~new_n3602_) & new_n3789_ & (~new_n3622_ | ~new_n3734_) & (new_n3718_ | ~P3_INSTQUEUE_REG_9__5__SCAN_IN);
  assign new_n3789_ = (~new_n3689_ | ~new_n3592_ | ~BUF2_REG_5__SCAN_IN) & (~new_n3627_ | ~BUF2_REG_21__SCAN_IN | ~new_n3592_ | ~new_n3725_);
  assign new_n3790_ = new_n3791_ & (~new_n2809_ | ~new_n2833_ | ~new_n2815_ | ~new_n2821_);
  assign new_n3791_ = new_n3602_ & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3792_ = (~new_n3624_ | new_n2833_ | ~new_n3602_) & new_n3795_ & ~new_n3794_ & (new_n3793_ | ~P3_INSTQUEUE_REG_13__4__SCAN_IN);
  assign new_n3793_ = ((~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) | (new_n3720_ & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)) & new_n3592_ & (~P3_STATE2_REG_3__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN));
  assign new_n3794_ = new_n3599_ & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & (~new_n3720_ | (new_n3725_ & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)));
  assign new_n3795_ = (~new_n3600_ | ~new_n3739_) & (~new_n3601_ | ~new_n3614_);
  assign new_n3796_ = new_n3797_ & (new_n3799_ | ~P3_INSTQUEUE_REG_5__0__SCAN_IN) & (~new_n3631_ | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  assign new_n3797_ = (~new_n3748_ | ~new_n3617_) & (~new_n3798_ | new_n3593_ | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  assign new_n3798_ = BUF2_REG_0__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & ((P3_STATE2_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (P3_STATE2_REG_2__SCAN_IN ^ P3_STATE2_REG_1__SCAN_IN));
  assign new_n3799_ = ((~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) | (new_n3720_ & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)) & new_n3592_ & (~P3_STATE2_REG_3__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN));
  assign new_n3800_ = new_n3803_ & ~new_n3801_ & ((P2_DATAO_REG_5__SCAN_IN & ~new_n3604_ & new_n3606_) | (new_n3604_ & P1_DATAO_REG_5__SCAN_IN) | (BUF1_REG_5__SCAN_IN & ~new_n3604_ & ~new_n3606_));
  assign new_n3801_ = new_n3802_ & (new_n3746_ | ~P3_INSTQUEUE_REG_2__0__SCAN_IN) & (~new_n3748_ | new_n2809_ | ~new_n3602_);
  assign new_n3802_ = (~new_n3631_ | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (~new_n3617_ | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (~new_n3798_ | new_n3593_ | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN));
  assign new_n3803_ = (new_n3804_ | ~new_n3805_ | (new_n3632_ & ~new_n2809_ & new_n3602_)) & (~new_n3748_ | ((new_n2815_ | ~new_n3602_) & (new_n2826_ | ~new_n3602_)));
  assign new_n3804_ = P3_INSTQUEUE_REG_4__0__SCAN_IN & (((P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) | (~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & (~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))) & (~new_n3720_ | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))) | ~new_n3592_ | (P3_STATE2_REG_3__SCAN_IN & (P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN)));
  assign new_n3805_ = (~new_n3629_ | ~new_n3798_) & (~new_n3617_ | ~new_n3692_) & (~new_n3748_ | ~new_n3631_);
  assign new_n3806_ = ~new_n3807_ & ~new_n3809_ & ((P2_DATAO_REG_0__SCAN_IN & ~new_n3604_ & new_n3606_) | (new_n3604_ & P1_DATAO_REG_0__SCAN_IN) | (BUF1_REG_0__SCAN_IN & ~new_n3604_ & ~new_n3606_));
  assign new_n3807_ = new_n3808_ & (new_n3736_ | ~P3_INSTQUEUE_REG_10__3__SCAN_IN) & (~new_n3739_ | new_n2821_ | ~new_n3602_);
  assign new_n3808_ = (~new_n3740_ | ~new_n3592_ | ~BUF2_REG_3__SCAN_IN) & (~new_n3620_ | ~BUF2_REG_19__SCAN_IN | ~new_n3592_ | ~new_n3725_) & (~new_n3627_ | ~BUF2_REG_27__SCAN_IN | ~new_n3592_ | ~new_n3725_);
  assign new_n3809_ = (~new_n3604_ | ~P1_DATAO_REG_3__SCAN_IN) & (~BUF1_REG_3__SCAN_IN | new_n3604_ | new_n3606_) & (~P2_DATAO_REG_3__SCAN_IN | new_n3604_ | ~new_n3606_);
  assign new_n3810_ = new_n3816_ & (~new_n3811_ | (new_n3614_ & ~new_n2826_ & new_n3602_)) & (~new_n3813_ | (new_n3733_ & ~new_n2796_ & new_n3602_));
  assign new_n3811_ = (new_n3783_ | ~P3_INSTQUEUE_REG_11__7__SCAN_IN) & (~new_n3616_ | ~new_n3620_) & ~new_n3812_ & (~new_n3628_ | ~new_n3630_);
  assign new_n3812_ = new_n3705_ & new_n3592_ & BUF2_REG_7__SCAN_IN;
  assign new_n3813_ = new_n3814_ & ~new_n3815_ & (new_n3799_ | ~P3_INSTQUEUE_REG_5__5__SCAN_IN);
  assign new_n3814_ = (~new_n3622_ | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (~new_n3592_ | ~BUF2_REG_5__SCAN_IN | new_n3593_ | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  assign new_n3815_ = new_n3591_ & BUF2_REG_21__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign new_n3816_ = (new_n3817_ | ~new_n3818_ | (~new_n3783_ & P3_INSTQUEUE_REG_11__2__SCAN_IN)) & (new_n3819_ | ~new_n3820_ | ~new_n3821_);
  assign new_n3817_ = new_n3614_ & new_n3602_ & (~new_n2816_ | ~new_n2817_ | ~new_n2818_ | ~new_n2819_ | ~new_n2820_);
  assign new_n3818_ = (~new_n3620_ | ~new_n3591_ | ~BUF2_REG_26__SCAN_IN) & (~new_n3738_ | ~new_n3705_) & (~new_n3630_ | ~new_n3591_ | ~BUF2_REG_18__SCAN_IN);
  assign new_n3819_ = new_n3630_ & new_n3602_ & (~new_n2834_ | ~new_n2835_ | ~new_n2836_ | ~new_n2837_ | ~new_n2838_);
  assign new_n3820_ = (~new_n3627_ | ~new_n3601_) & (~new_n3599_ | ~new_n3689_);
  assign new_n3821_ = (~new_n3600_ | ~new_n3734_) & (~P3_INSTQUEUE_REG_9__4__SCAN_IN | (new_n3592_ & ~new_n3621_));
  assign new_n3822_ = ~new_n3823_ & ~new_n3825_ & ~new_n3828_ & (new_n3824_ | new_n3581_ | ~new_n2950_);
  assign new_n3823_ = (~new_n3585_ | new_n1322_ | (new_n2976_ ? ~BUF1_REG_1__SCAN_IN : ~BUF2_REG_1__SCAN_IN)) & (~new_n3440_ | ~P2_EAX_REG_17__SCAN_IN) & (new_n3585_ | ~P2_UWORD_REG_1__SCAN_IN);
  assign new_n3824_ = (new_n2945_ | (~new_n2928_ & ~new_n2850_)) & (new_n3582_ | new_n3446_) & (~new_n2927_ | new_n2939_);
  assign new_n3825_ = ~new_n3827_ & (~new_n2950_ | (~new_n3826_ & (~new_n2854_ | ~new_n2945_)));
  assign new_n3826_ = ~new_n2802_ & ~new_n2809_ & new_n2826_ & new_n2833_ & new_n2815_ & new_n2821_ & ~new_n2790_ & new_n2796_;
  assign new_n3827_ = ~P3_EBX_REG_15__SCAN_IN & ~P3_EBX_REG_16__SCAN_IN & ~P3_EBX_REG_31__SCAN_IN & P3_EBX_REG_20__SCAN_IN & P3_EBX_REG_28__SCAN_IN;
  assign new_n3828_ = (~new_n3445_ | ((~new_n2839_ | ~new_n2802_) & (new_n2943_ | ~new_n2839_ | new_n2802_))) & (~new_n3829_ | P3_UWORD_REG_2__SCAN_IN | P3_UWORD_REG_13__SCAN_IN | P3_UWORD_REG_6__SCAN_IN);
  assign new_n3829_ = ~P3_LWORD_REG_9__SCAN_IN & ~P3_LWORD_REG_6__SCAN_IN & ~P3_LWORD_REG_3__SCAN_IN & ~P3_LWORD_REG_1__SCAN_IN & ~P3_LWORD_REG_14__SCAN_IN & ~P3_LWORD_REG_13__SCAN_IN & ~P3_LWORD_REG_10__SCAN_IN & ~P3_UWORD_REG_9__SCAN_IN;
  assign new_n3830_ = ~new_n3836_ & ~new_n3882_ & ~new_n3831_ & ~new_n3832_ & ~new_n3883_ & ~new_n3885_ & ~new_n3886_ & ~new_n3887_;
  assign new_n3831_ = (~P3_UWORD_REG_1__SCAN_IN | (new_n3445_ & ((new_n2839_ & new_n2802_) | ((~READY2 | ~READY22_REG_SCAN_IN) & new_n2839_ & ~new_n2802_)))) & (~BUF2_REG_1__SCAN_IN | ~new_n3445_ | (READY2 & READY22_REG_SCAN_IN) | ~new_n2839_ | new_n2802_) & (~P3_EAX_REG_17__SCAN_IN | ~new_n3445_ | ~new_n2839_ | ~new_n2802_);
  assign new_n3832_ = new_n2826_ & new_n2950_ & (new_n3826_ | (new_n2854_ & new_n2945_)) & (~new_n3833_ | ~P3_EBX_REG_15__SCAN_IN | ~P3_EBX_REG_16__SCAN_IN) & ((new_n3833_ & P3_EBX_REG_15__SCAN_IN) | P3_EBX_REG_16__SCAN_IN);
  assign new_n3833_ = new_n3834_ & new_n3835_;
  assign new_n3834_ = P3_EBX_REG_5__SCAN_IN & P3_EBX_REG_6__SCAN_IN & P3_EBX_REG_3__SCAN_IN & P3_EBX_REG_4__SCAN_IN & P3_EBX_REG_7__SCAN_IN & P3_EBX_REG_8__SCAN_IN & P3_EBX_REG_9__SCAN_IN & P3_EBX_REG_10__SCAN_IN;
  assign new_n3835_ = P3_EBX_REG_2__SCAN_IN & P3_EBX_REG_0__SCAN_IN & P3_EBX_REG_1__SCAN_IN & P3_EBX_REG_13__SCAN_IN & P3_EBX_REG_14__SCAN_IN & P3_EBX_REG_11__SCAN_IN & P3_EBX_REG_12__SCAN_IN;
  assign new_n3836_ = (new_n3837_ | new_n2826_ | new_n3877_) & ~new_n3873_ & new_n2950_ & (new_n3826_ | (new_n2854_ & new_n2945_));
  assign new_n3837_ = new_n3868_ ^ (~new_n3858_ & ~new_n3863_ & ~new_n3853_ & ~new_n3848_ & ~new_n3838_ & ~new_n3843_);
  assign new_n3838_ = new_n3840_ & new_n3841_ & new_n3842_ & new_n3839_ & (~new_n2868_ | ~P3_INSTQUEUE_REG_1__7__SCAN_IN) & (~new_n2804_ | ~P3_INSTQUEUE_REG_2__7__SCAN_IN);
  assign new_n3839_ = (~P3_INSTQUEUE_REG_10__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_14__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_3__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3840_ = (~P3_INSTQUEUE_REG_9__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_11__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3841_ = (~P3_INSTQUEUE_REG_7__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_8__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3842_ = (~P3_INSTQUEUE_REG_12__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_0__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_5__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_15__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3843_ = new_n3845_ & new_n3846_ & new_n3847_ & new_n3844_ & (~new_n2868_ | ~P3_INSTQUEUE_REG_2__0__SCAN_IN) & (~new_n2803_ | ~P3_INSTQUEUE_REG_11__0__SCAN_IN);
  assign new_n3844_ = (~P3_INSTQUEUE_REG_3__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_15__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3845_ = (~P3_INSTQUEUE_REG_10__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_5__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3846_ = (~P3_INSTQUEUE_REG_0__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_4__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_1__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_7__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3847_ = (~P3_INSTQUEUE_REG_12__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_14__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_8__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3848_ = new_n3850_ & new_n3851_ & new_n3852_ & new_n3849_ & (~new_n2804_ | ~P3_INSTQUEUE_REG_3__1__SCAN_IN) & (~new_n2803_ | ~P3_INSTQUEUE_REG_11__1__SCAN_IN);
  assign new_n3849_ = (~P3_INSTQUEUE_REG_2__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_4__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_7__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3850_ = (~P3_INSTQUEUE_REG_0__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_12__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3851_ = (~P3_INSTQUEUE_REG_10__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3852_ = (~P3_INSTQUEUE_REG_5__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_15__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_14__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_1__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3853_ = new_n3855_ & new_n3856_ & new_n3857_ & new_n3854_ & (~new_n2868_ | ~P3_INSTQUEUE_REG_2__2__SCAN_IN) & (~new_n2803_ | ~P3_INSTQUEUE_REG_11__2__SCAN_IN);
  assign new_n3854_ = (~P3_INSTQUEUE_REG_3__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_4__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3855_ = (~P3_INSTQUEUE_REG_10__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_5__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3856_ = (~P3_INSTQUEUE_REG_8__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_0__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_7__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_1__2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3857_ = (~P3_INSTQUEUE_REG_15__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_14__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3858_ = new_n3860_ & new_n3861_ & new_n3862_ & new_n3859_ & (~new_n2868_ | ~P3_INSTQUEUE_REG_2__3__SCAN_IN) & (~new_n2804_ | ~P3_INSTQUEUE_REG_3__3__SCAN_IN);
  assign new_n3859_ = (~P3_INSTQUEUE_REG_11__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_15__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3860_ = (~P3_INSTQUEUE_REG_0__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_8__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3861_ = (~P3_INSTQUEUE_REG_10__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_5__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_1__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3862_ = (~P3_INSTQUEUE_REG_12__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_14__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_7__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3863_ = new_n3865_ & new_n3866_ & new_n3867_ & new_n3864_ & (~new_n2804_ | ~P3_INSTQUEUE_REG_3__4__SCAN_IN) & (~new_n2803_ | ~P3_INSTQUEUE_REG_11__4__SCAN_IN);
  assign new_n3864_ = (~P3_INSTQUEUE_REG_2__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_6__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3865_ = (~P3_INSTQUEUE_REG_0__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_10__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3866_ = (~P3_INSTQUEUE_REG_5__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_15__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_14__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_1__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3867_ = (~P3_INSTQUEUE_REG_9__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_7__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_12__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_4__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3868_ = new_n3870_ & new_n3871_ & new_n3872_ & new_n3869_ & (~new_n2868_ | ~P3_INSTQUEUE_REG_2__5__SCAN_IN) & (~new_n2803_ | ~P3_INSTQUEUE_REG_11__5__SCAN_IN);
  assign new_n3869_ = (~P3_INSTQUEUE_REG_3__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_4__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_5__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3870_ = (~P3_INSTQUEUE_REG_15__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_6__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3871_ = (~P3_INSTQUEUE_REG_8__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_1__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_14__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3872_ = (~P3_INSTQUEUE_REG_10__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_0__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_7__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3873_ = (~P3_EBX_REG_28__SCAN_IN | ~new_n3876_ | ~P3_EBX_REG_21__SCAN_IN | ~new_n3874_ | ~P3_EBX_REG_20__SCAN_IN) & (P3_EBX_REG_28__SCAN_IN | (new_n3876_ & P3_EBX_REG_21__SCAN_IN & new_n3874_ & P3_EBX_REG_20__SCAN_IN)) & (new_n3874_ | P3_EBX_REG_20__SCAN_IN) & new_n2826_ & (~new_n3874_ | ~P3_EBX_REG_20__SCAN_IN);
  assign new_n3874_ = new_n3875_ & P3_EBX_REG_17__SCAN_IN & P3_EBX_REG_16__SCAN_IN & P3_EBX_REG_15__SCAN_IN & new_n3834_ & new_n3835_;
  assign new_n3875_ = P3_EBX_REG_18__SCAN_IN & P3_EBX_REG_19__SCAN_IN;
  assign new_n3876_ = P3_EBX_REG_22__SCAN_IN & P3_EBX_REG_25__SCAN_IN & P3_EBX_REG_26__SCAN_IN & P3_EBX_REG_27__SCAN_IN & P3_EBX_REG_23__SCAN_IN & P3_EBX_REG_24__SCAN_IN;
  assign new_n3877_ = new_n3879_ & new_n3880_ & new_n3881_ & new_n3878_ & (~new_n2868_ | ~P3_INSTQUEUE_REG_1__4__SCAN_IN) & (~new_n2804_ | ~P3_INSTQUEUE_REG_2__4__SCAN_IN);
  assign new_n3878_ = (~P3_INSTQUEUE_REG_10__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3879_ = (~P3_INSTQUEUE_REG_11__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_14__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3880_ = (~P3_INSTQUEUE_REG_7__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_3__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_15__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3881_ = (~P3_INSTQUEUE_REG_6__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_0__4__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_13__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_5__4__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3882_ = new_n3585_ & ~new_n1322_ & (new_n2976_ | BUF2_REG_15__SCAN_IN) & (~new_n2976_ | BUF1_REG_15__SCAN_IN);
  assign new_n3883_ = ~new_n3884_ & new_n3448_ & (~new_n3445_ | new_n3447_);
  assign new_n3884_ = ~P3_REIP_REG_25__SCAN_IN & ~P3_REIP_REG_30__SCAN_IN & ~P3_REIP_REG_7__SCAN_IN & ~P3_REIP_REG_10__SCAN_IN & ~P3_REIP_REG_1__SCAN_IN & ~P3_REIP_REG_3__SCAN_IN;
  assign new_n3885_ = (~P3_UWORD_REG_12__SCAN_IN | (new_n3445_ & ((new_n2839_ & new_n2802_) | ((~READY2 | ~READY22_REG_SCAN_IN) & new_n2839_ & ~new_n2802_)))) & (~BUF2_REG_12__SCAN_IN | ~new_n3445_ | (READY2 & READY22_REG_SCAN_IN) | ~new_n2839_ | new_n2802_) & (~P3_EAX_REG_28__SCAN_IN | ~new_n3445_ | ~new_n2839_ | ~new_n2802_);
  assign new_n3886_ = (~P3_UWORD_REG_10__SCAN_IN | (new_n3445_ & ((new_n2839_ & new_n2802_) | ((~READY2 | ~READY22_REG_SCAN_IN) & new_n2839_ & ~new_n2802_)))) & (~BUF2_REG_10__SCAN_IN | ~new_n3445_ | (READY2 & READY22_REG_SCAN_IN) | ~new_n2839_ | new_n2802_) & (~P3_EAX_REG_26__SCAN_IN | ~new_n3445_ | ~new_n2839_ | ~new_n2802_);
  assign new_n3887_ = (~P3_LWORD_REG_8__SCAN_IN | (new_n3445_ & ((new_n2839_ & new_n2802_) | ((~READY2 | ~READY22_REG_SCAN_IN) & new_n2839_ & ~new_n2802_)))) & (~BUF2_REG_8__SCAN_IN | ~new_n3445_ | (READY2 & READY22_REG_SCAN_IN) | ~new_n2839_ | new_n2802_) & (~P3_EAX_REG_8__SCAN_IN | ~new_n3445_ | ~new_n2839_ | ~new_n2802_);
  assign new_n3888_ = ~new_n3891_ & ~new_n3892_ & ~new_n3890_ & (~new_n3889_ | (~P3_LWORD_REG_10__SCAN_IN & ~P3_UWORD_REG_9__SCAN_IN & ~P3_UWORD_REG_5__SCAN_IN & ~P3_UWORD_REG_2__SCAN_IN));
  assign new_n3889_ = ~P3_STATE2_REG_0__SCAN_IN & ((new_n3445_ & new_n2947_ & (new_n2840_ | new_n3518_)) | (P3_STATE2_REG_1__SCAN_IN & P3_STATE2_REG_2__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN));
  assign new_n3890_ = (~new_n3585_ | new_n1322_ | (new_n2976_ ? ~BUF1_REG_10__SCAN_IN : ~BUF2_REG_10__SCAN_IN)) & (~new_n3440_ | ~P2_EAX_REG_10__SCAN_IN) & (new_n3585_ | ~P2_LWORD_REG_10__SCAN_IN);
  assign new_n3891_ = (~new_n3585_ | new_n1322_ | (new_n2976_ ? ~BUF1_REG_7__SCAN_IN : ~BUF2_REG_7__SCAN_IN)) & (~new_n3440_ | ~P2_EAX_REG_23__SCAN_IN) & (new_n3585_ | ~P2_UWORD_REG_7__SCAN_IN);
  assign new_n3892_ = (new_n3893_ | ~new_n2950_ | (~new_n3826_ & (~new_n2854_ | ~new_n2945_))) & (~P3_EBX_REG_22__SCAN_IN | ~P3_EBX_REG_25__SCAN_IN | (~new_n3901_ & new_n2950_ & (new_n3826_ | (new_n2854_ & new_n2945_))));
  assign new_n3893_ = ((new_n3853_ & (new_n3848_ | new_n3838_ | new_n3843_)) | new_n2826_ | new_n3895_ | (~new_n3853_ & ~new_n3848_ & ~new_n3838_ & ~new_n3843_)) & (~new_n3894_ | ~new_n2826_ | ~new_n3900_);
  assign new_n3894_ = P3_EBX_REG_21__SCAN_IN & P3_EBX_REG_20__SCAN_IN & new_n3875_ & P3_EBX_REG_17__SCAN_IN & P3_EBX_REG_16__SCAN_IN & P3_EBX_REG_15__SCAN_IN & new_n3834_ & new_n3835_;
  assign new_n3895_ = new_n3897_ & new_n3898_ & new_n3899_ & new_n3896_ & (~new_n2868_ | ~P3_INSTQUEUE_REG_1__6__SCAN_IN) & (~new_n2804_ | ~P3_INSTQUEUE_REG_2__6__SCAN_IN);
  assign new_n3896_ = (~P3_INSTQUEUE_REG_10__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3897_ = (~P3_INSTQUEUE_REG_11__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_14__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3898_ = (~P3_INSTQUEUE_REG_7__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_3__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_15__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3899_ = (~P3_INSTQUEUE_REG_6__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_0__6__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_13__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_5__6__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3900_ = ~P3_EBX_REG_22__SCAN_IN & P3_EBX_REG_25__SCAN_IN;
  assign new_n3901_ = new_n2826_ & ~new_n3894_;
  assign new_n3902_ = ~new_n3905_ & ~new_n3906_ & ~new_n3903_ & ~new_n3904_;
  assign new_n3903_ = (~new_n3585_ | new_n1322_ | (new_n2976_ ? ~BUF1_REG_3__SCAN_IN : ~BUF2_REG_3__SCAN_IN)) & (~new_n3440_ | ~P2_EAX_REG_19__SCAN_IN) & (new_n3585_ | ~P2_UWORD_REG_3__SCAN_IN);
  assign new_n3904_ = (~new_n3585_ | new_n1322_ | (new_n2976_ ? ~BUF1_REG_0__SCAN_IN : ~BUF2_REG_0__SCAN_IN)) & (~new_n3440_ | ~P2_EAX_REG_0__SCAN_IN) & (new_n3585_ | ~P2_LWORD_REG_0__SCAN_IN);
  assign new_n3905_ = (new_n3585_ | ~P2_UWORD_REG_5__SCAN_IN) & (~new_n3440_ | ~P2_EAX_REG_21__SCAN_IN) & (new_n3078_ | ~new_n3585_ | new_n1322_);
  assign new_n3906_ = (~new_n3585_ | new_n1322_ | (new_n2976_ ? ~BUF1_REG_2__SCAN_IN : ~BUF2_REG_2__SCAN_IN)) & (~new_n3440_ | ~P2_EAX_REG_2__SCAN_IN) & (new_n3585_ | ~P2_LWORD_REG_2__SCAN_IN);
  assign new_n3907_ = new_n3908_ & ~new_n3917_ & (~new_n3516_ | ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) & ~new_n3920_ & (new_n3516_ | ~new_n3923_ | ~new_n2832_ | (new_n3921_ & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (~new_n3921_ & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN));
  assign new_n3908_ = ~new_n3909_ & (~BUF2_REG_21__SCAN_IN | ~new_n3912_ | new_n2790_) & ~new_n3913_ & (~BUF2_REG_5__SCAN_IN | ~new_n3912_ | (new_n2790_ & ~new_n2796_));
  assign new_n3909_ = ~new_n3911_ & new_n3910_ & new_n3472_ & P3_STATE2_REG_2__SCAN_IN & (~new_n3448_ | (new_n3445_ & ~new_n3447_));
  assign new_n3910_ = new_n3474_ & new_n2947_;
  assign new_n3911_ = P3_REIP_REG_1__SCAN_IN & (~new_n3485_ ^ P3_REIP_REG_25__SCAN_IN) & (~P3_REIP_REG_3__SCAN_IN ^ (P3_REIP_REG_1__SCAN_IN & P3_REIP_REG_2__SCAN_IN));
  assign new_n3912_ = ~new_n2826_ & new_n2950_ & (new_n3525_ | (new_n2853_ & new_n2945_) | (~new_n3520_ & new_n2942_));
  assign new_n3913_ = ~new_n3914_ & new_n3474_ & new_n3473_ & P3_STATE2_REG_2__SCAN_IN & (~new_n3448_ | (new_n3445_ & ~new_n3447_));
  assign new_n3914_ = new_n3915_ & (~P3_REIP_REG_3__SCAN_IN ^ (P3_REIP_REG_1__SCAN_IN & P3_REIP_REG_2__SCAN_IN)) & (~new_n3485_ ^ P3_REIP_REG_25__SCAN_IN);
  assign new_n3915_ = (~new_n3916_ ^ P3_REIP_REG_7__SCAN_IN) & (~P3_REIP_REG_10__SCAN_IN ^ (P3_REIP_REG_9__SCAN_IN & P3_REIP_REG_8__SCAN_IN & new_n3916_ & P3_REIP_REG_7__SCAN_IN));
  assign new_n3916_ = P3_REIP_REG_3__SCAN_IN & P3_REIP_REG_1__SCAN_IN & P3_REIP_REG_2__SCAN_IN & P3_REIP_REG_6__SCAN_IN & P3_REIP_REG_4__SCAN_IN & P3_REIP_REG_5__SCAN_IN;
  assign new_n3917_ = (~P3_INSTQUEUE_REG_0__4__SCAN_IN | ~new_n3918_ | new_n2826_) & ((P3_EBX_REG_4__SCAN_IN & new_n3918_ & new_n3919_ & P3_EBX_REG_3__SCAN_IN) | (new_n3918_ & ~new_n2826_) | (~P3_EBX_REG_4__SCAN_IN & (~new_n3918_ | ~new_n3919_ | ~P3_EBX_REG_3__SCAN_IN)));
  assign new_n3918_ = new_n2950_ & (new_n3826_ | (new_n2854_ & new_n2945_));
  assign new_n3919_ = P3_EBX_REG_2__SCAN_IN & P3_EBX_REG_0__SCAN_IN & P3_EBX_REG_1__SCAN_IN;
  assign new_n3920_ = BUF2_REG_8__SCAN_IN & new_n3912_ & ~new_n3522_;
  assign new_n3921_ = new_n3922_ & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign new_n3922_ = P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign new_n3923_ = ~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_1__SCAN_IN;
  assign new_n3924_ = ~new_n3925_ & (new_n3935_ | new_n2937_ | new_n3282_) & (new_n3929_ | ~new_n2937_) & (~new_n2005_ | (~P2_PHYADDRPOINTER_REG_13__SCAN_IN & ~P2_PHYADDRPOINTER_REG_17__SCAN_IN));
  assign new_n3925_ = (new_n3296_ | P3_PHYADDRPOINTER_REG_1__SCAN_IN) & (~P3_PHYADDRPOINTER_REG_1__SCAN_IN | (~new_n3293_ & ~new_n3305_)) & new_n3926_ & (~P3_REIP_REG_1__SCAN_IN | new_n3293_ | ~new_n3284_);
  assign new_n3926_ = (new_n3927_ | ~new_n2802_ | ~new_n2950_ | ((~new_n2927_ | ~new_n2939_) & (~new_n2928_ | ~new_n2945_))) & (new_n3928_ | new_n2802_ | ~new_n2950_ | ((~new_n2927_ | ~new_n2939_) & (~new_n2928_ | ~new_n2945_)));
  assign new_n3927_ = (~new_n2883_ | P3_INSTADDRPOINTER_REG_0__SCAN_IN) ^ (new_n2873_ ^ P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  assign new_n3928_ = ~new_n2919_ ^ (new_n2873_ ^ P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  assign new_n3929_ = (new_n3286_ | (new_n2844_ & P3_INSTADDRPOINTER_REG_3__SCAN_IN) | (~new_n2844_ & ~P3_INSTADDRPOINTER_REG_3__SCAN_IN)) & new_n3930_ & ((~new_n3934_ & (P3_INSTADDRPOINTER_REG_3__SCAN_IN ^ (~new_n3933_ ^ new_n2878_))) | ~new_n2928_ | (new_n3934_ & (P3_INSTADDRPOINTER_REG_3__SCAN_IN | (new_n3933_ ^ new_n2878_)) & (~P3_INSTADDRPOINTER_REG_3__SCAN_IN | (new_n3933_ & new_n2878_) | (~new_n3933_ & ~new_n2878_))));
  assign new_n3930_ = ((new_n3932_ & (new_n3931_ | P3_INSTADDRPOINTER_REG_3__SCAN_IN) & (~new_n3931_ | ~P3_INSTADDRPOINTER_REG_3__SCAN_IN)) | ~new_n2927_ | (~new_n3932_ & (new_n3931_ ^ ~P3_INSTADDRPOINTER_REG_3__SCAN_IN))) & (~new_n2850_ | (new_n2849_ & ~P3_INSTADDRPOINTER_REG_3__SCAN_IN) | (~new_n2849_ & P3_INSTADDRPOINTER_REG_3__SCAN_IN)) & (new_n3287_ | (new_n2785_ & P3_INSTADDRPOINTER_REG_3__SCAN_IN) | (~new_n2785_ & ~P3_INSTADDRPOINTER_REG_3__SCAN_IN));
  assign new_n3931_ = ~new_n2878_ ^ (~new_n2867_ & ~new_n2873_);
  assign new_n3932_ = (P3_INSTADDRPOINTER_REG_2__SCAN_IN | (new_n2867_ ^ new_n2873_)) & ((P3_INSTADDRPOINTER_REG_2__SCAN_IN & (~new_n2867_ | ~new_n2873_) & (new_n2867_ | new_n2873_)) | ((new_n2919_ | (new_n2873_ & P3_INSTADDRPOINTER_REG_1__SCAN_IN)) & (new_n2873_ | P3_INSTADDRPOINTER_REG_1__SCAN_IN)));
  assign new_n3933_ = new_n2867_ & (new_n2873_ | new_n2883_);
  assign new_n3934_ = (P3_INSTADDRPOINTER_REG_2__SCAN_IN | (~new_n2867_ & ~new_n2873_ & ~new_n2883_) | (new_n2867_ & (new_n2873_ | new_n2883_))) & ((P3_INSTADDRPOINTER_REG_2__SCAN_IN & (new_n2867_ ^ (~new_n2873_ & ~new_n2883_))) | (((~new_n2873_ & P3_INSTADDRPOINTER_REG_1__SCAN_IN) | ~new_n2883_ | P3_INSTADDRPOINTER_REG_0__SCAN_IN) & (new_n2873_ | new_n2883_) & (~new_n2873_ | P3_INSTADDRPOINTER_REG_1__SCAN_IN)));
  assign new_n3935_ = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN & ~P3_INSTADDRPOINTER_REG_31__SCAN_IN & ~P3_INSTADDRPOINTER_REG_25__SCAN_IN & ~P3_INSTADDRPOINTER_REG_3__SCAN_IN & ~P3_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign new_n3936_ = ~new_n3978_ & new_n3983_ & new_n3985_ & new_n3937_ & new_n3975_ & new_n3956_ & new_n3966_ & new_n3973_;
  assign new_n3937_ = ~new_n3948_ & ~new_n3955_ & (new_n3296_ | ~new_n3459_) & (new_n3938_ | ~new_n3565_ | ~new_n3522_);
  assign new_n3938_ = new_n3837_ & (new_n3838_ ^ ~new_n3843_) & new_n2894_ & new_n3939_ & new_n3945_ & new_n3946_ & new_n3947_;
  assign new_n3939_ = new_n3941_ & new_n3943_ & new_n3944_ & new_n3940_ & (~new_n2803_ | (~P3_INSTQUEUE_REG_10__5__SCAN_IN & ~P3_INSTQUEUE_REG_9__0__SCAN_IN));
  assign new_n3940_ = (~new_n2804_ | ~P3_INSTQUEUE_REG_1__0__SCAN_IN) & (~new_n2868_ | (~P3_INSTQUEUE_REG_1__5__SCAN_IN & ~P3_INSTQUEUE_REG_0__0__SCAN_IN));
  assign new_n3941_ = new_n3942_ & (~P3_INSTQUEUE_REG_2__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_8__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_0__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3942_ = (~P3_INSTQUEUE_REG_13__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_4__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_6__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3943_ = (~P3_INSTQUEUE_REG_2__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_4__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_7__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_11__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3944_ = (~P3_INSTQUEUE_REG_8__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_5__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_10__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_3__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3945_ = (~P3_INSTQUEUE_REG_7__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_14__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_14__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3946_ = (~P3_INSTQUEUE_REG_13__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_15__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_11__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3947_ = (~P3_INSTQUEUE_REG_5__5__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_15__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_3__5__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3948_ = (~new_n2826_ | ~new_n2950_ | (~new_n3826_ & (~new_n2854_ | ~new_n2945_)) | (new_n3949_ & P3_EBX_REG_17__SCAN_IN) | (~new_n3949_ & ~P3_EBX_REG_17__SCAN_IN)) & (new_n3950_ | new_n2826_ | ~new_n2950_ | (~new_n3826_ & (~new_n2854_ | ~new_n2945_))) & (~P3_EBX_REG_17__SCAN_IN | (new_n2950_ & (new_n3826_ | (new_n2854_ & new_n2945_))));
  assign new_n3949_ = P3_EBX_REG_16__SCAN_IN & new_n3833_ & P3_EBX_REG_15__SCAN_IN;
  assign new_n3950_ = new_n3952_ & new_n3953_ & new_n3954_ & new_n3951_ & (~new_n2868_ | ~P3_INSTQUEUE_REG_1__1__SCAN_IN) & (~new_n2804_ | ~P3_INSTQUEUE_REG_2__1__SCAN_IN);
  assign new_n3951_ = (~P3_INSTQUEUE_REG_10__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3952_ = (~P3_INSTQUEUE_REG_11__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_14__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3953_ = (~P3_INSTQUEUE_REG_7__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_12__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_3__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_15__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3954_ = (~P3_INSTQUEUE_REG_6__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_0__1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_13__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_5__1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3955_ = ((new_n3919_ & P3_EBX_REG_3__SCAN_IN) | (~new_n3919_ & ~P3_EBX_REG_3__SCAN_IN) | ~new_n2826_ | ~new_n2950_ | (~new_n3826_ & (~new_n2854_ | ~new_n2945_))) & (~P3_INSTQUEUE_REG_0__3__SCAN_IN | new_n2826_ | ~new_n2950_ | (~new_n3826_ & (~new_n2854_ | ~new_n2945_))) & (~P3_EBX_REG_3__SCAN_IN | (new_n2950_ & (new_n3826_ | (new_n2854_ & new_n2945_))));
  assign new_n3956_ = ~new_n3959_ & (~new_n3957_ | (new_n3833_ & P3_EBX_REG_15__SCAN_IN) | (~new_n3833_ & ~P3_EBX_REG_15__SCAN_IN)) & (~new_n3293_ | new_n3965_) & (~new_n3958_ | new_n3960_);
  assign new_n3957_ = new_n2826_ & new_n2950_ & (new_n3826_ | (new_n2854_ & new_n2945_));
  assign new_n3958_ = ~new_n2826_ & new_n2950_ & (new_n3826_ | (new_n2854_ & new_n2945_));
  assign new_n3959_ = (~P3_UWORD_REG_14__SCAN_IN | (new_n3445_ & ((new_n2839_ & new_n2802_) | ((~READY2 | ~READY22_REG_SCAN_IN) & new_n2839_ & ~new_n2802_)))) & (~BUF2_REG_14__SCAN_IN | ~new_n3445_ | (READY2 & READY22_REG_SCAN_IN) | ~new_n2839_ | new_n2802_) & (~P3_EAX_REG_30__SCAN_IN | ~new_n3445_ | ~new_n2839_ | ~new_n2802_);
  assign new_n3960_ = new_n3962_ & new_n3963_ & new_n3964_ & new_n3961_ & (~new_n2868_ | ~P3_INSTQUEUE_REG_0__7__SCAN_IN) & (~new_n2803_ | ~P3_INSTQUEUE_REG_9__7__SCAN_IN);
  assign new_n3961_ = (~P3_INSTQUEUE_REG_1__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_15__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_3__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3962_ = (~P3_INSTQUEUE_REG_4__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_12__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3963_ = (~P3_INSTQUEUE_REG_11__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_8__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_7__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3964_ = (~P3_INSTQUEUE_REG_2__7__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_5__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_10__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_14__7__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3965_ = ~P3_PHYADDRPOINTER_REG_21__SCAN_IN & ~P3_PHYADDRPOINTER_REG_12__SCAN_IN & ~P3_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign new_n3966_ = (~new_n3958_ | new_n3968_) & (~new_n3967_ | (~P3_DATAO_REG_10__SCAN_IN & ~P3_DATAO_REG_18__SCAN_IN & ~P3_DATAO_REG_21__SCAN_IN & ~P3_DATAO_REG_25__SCAN_IN));
  assign new_n3967_ = (~new_n3297_ | ~P3_STATE2_REG_1__SCAN_IN) & (~new_n3445_ | ~new_n2947_ | (~new_n2840_ & ~new_n3518_));
  assign new_n3968_ = new_n3970_ & new_n3971_ & new_n3972_ & new_n3969_ & (~new_n2868_ | ~P3_INSTQUEUE_REG_1__0__SCAN_IN) & (~new_n2804_ | ~P3_INSTQUEUE_REG_2__0__SCAN_IN);
  assign new_n3969_ = (~P3_INSTQUEUE_REG_10__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_7__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_8__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3970_ = (~P3_INSTQUEUE_REG_11__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_4__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_14__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3971_ = (~P3_INSTQUEUE_REG_5__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_15__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_6__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_0__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n3972_ = (~P3_INSTQUEUE_REG_12__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_3__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_9__0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_13__0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n3973_ = ~new_n3974_ & (~new_n3957_ | (~P3_EBX_REG_31__SCAN_IN & (~new_n3894_ | ~new_n3876_ | ~P3_EBX_REG_30__SCAN_IN | ~P3_EBX_REG_28__SCAN_IN | ~P3_EBX_REG_29__SCAN_IN)) | (P3_EBX_REG_31__SCAN_IN & new_n3894_ & new_n3876_ & P3_EBX_REG_30__SCAN_IN & P3_EBX_REG_28__SCAN_IN & P3_EBX_REG_29__SCAN_IN));
  assign new_n3974_ = (P3_EAX_REG_18__SCAN_IN | P3_EAX_REG_21__SCAN_IN) & ~new_n2809_ & new_n3445_ & new_n2947_ & (new_n2840_ | new_n3518_);
  assign new_n3975_ = ~new_n2006_ & (~new_n3332_ | ~new_n3977_) & (~new_n3293_ | ~P3_PHYADDRPOINTER_REG_0__SCAN_IN) & (~new_n3976_ | ~P3_EAX_REG_25__SCAN_IN) & (~new_n3306_ | new_n3977_);
  assign new_n3976_ = ~new_n2809_ & new_n3445_ & new_n2947_ & (new_n2840_ | new_n3518_);
  assign new_n3977_ = new_n2883_ ^ ~P3_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign new_n3978_ = new_n3476_ & ~new_n3979_;
  assign new_n3979_ = (~P3_EBX_REG_30__SCAN_IN | ~new_n3982_ | P3_EBX_REG_27__SCAN_IN | P3_EBX_REG_26__SCAN_IN | P3_EBX_REG_25__SCAN_IN | ~new_n3478_ | ~new_n3482_) & (P3_EBX_REG_30__SCAN_IN | (new_n3982_ & ~P3_EBX_REG_27__SCAN_IN & ~P3_EBX_REG_26__SCAN_IN & ~P3_EBX_REG_25__SCAN_IN & new_n3478_ & new_n3482_)) & new_n3980_ & (~P3_EBX_REG_25__SCAN_IN ^ (~new_n3478_ | ~new_n3482_));
  assign new_n3980_ = new_n3981_ & (P3_EBX_REG_10__SCAN_IN ^ (~P3_EBX_REG_9__SCAN_IN & new_n3480_ & ~P3_EBX_REG_8__SCAN_IN));
  assign new_n3981_ = (P3_EBX_REG_7__SCAN_IN ^ (~P3_EBX_REG_6__SCAN_IN & ~P3_EBX_REG_4__SCAN_IN & ~P3_EBX_REG_5__SCAN_IN & ~P3_EBX_REG_3__SCAN_IN & ~P3_EBX_REG_2__SCAN_IN & ~P3_EBX_REG_0__SCAN_IN & ~P3_EBX_REG_1__SCAN_IN)) & (~P3_EBX_REG_0__SCAN_IN ^ P3_EBX_REG_1__SCAN_IN) & (P3_EBX_REG_3__SCAN_IN ^ (~P3_EBX_REG_2__SCAN_IN & ~P3_EBX_REG_0__SCAN_IN & ~P3_EBX_REG_1__SCAN_IN));
  assign new_n3982_ = ~P3_EBX_REG_28__SCAN_IN & ~P3_EBX_REG_29__SCAN_IN;
  assign new_n3983_ = ((new_n3976_ & P3_EAX_REG_23__SCAN_IN) | (new_n3967_ & P3_DATAO_REG_23__SCAN_IN) | (P3_UWORD_REG_7__SCAN_IN & ~new_n3967_ & ~P3_STATE2_REG_0__SCAN_IN)) & (~new_n3984_ | (P3_LWORD_REG_1__SCAN_IN & ~new_n3967_ & ~P3_STATE2_REG_0__SCAN_IN));
  assign new_n3984_ = (~P3_EAX_REG_1__SCAN_IN | ~new_n3445_ | ~new_n2947_ | (~new_n2840_ & ~new_n3518_)) & (~P3_DATAO_REG_1__SCAN_IN | (new_n3297_ & P3_STATE2_REG_1__SCAN_IN) | (new_n3445_ & new_n2947_ & (new_n2840_ | new_n3518_)));
  assign new_n3985_ = (~new_n3912_ | ~new_n2796_ | ~BUF2_REG_12__SCAN_IN) & (~new_n3912_ | ((~new_n2796_ | ~BUF2_REG_7__SCAN_IN) & (new_n2790_ | ~BUF2_REG_23__SCAN_IN)));
  assign new_n3986_ = (~new_n3439_ & (~new_n1407_ | ~P2_STATE2_REG_1__SCAN_IN)) ? (~P2_DATAO_REG_20__SCAN_IN & ~P2_DATAO_REG_7__SCAN_IN & ~P2_DATAO_REG_10__SCAN_IN) : (~new_n1340_ | ~P2_EAX_REG_20__SCAN_IN);
  assign new_n3987_ = new_n3988_ & new_n3996_ & new_n4007_ & ~new_n4023_ & (new_n2724_ | ~new_n3374_);
  assign new_n3988_ = new_n3989_ & ~new_n3993_ & (~new_n3509_ | (~P1_EAX_REG_7__SCAN_IN & ~P1_EAX_REG_15__SCAN_IN & ~P1_EAX_REG_14__SCAN_IN));
  assign new_n3989_ = (new_n3990_ | new_n3449_ | new_n3444_ | ~P3_STATE2_REG_1__SCAN_IN) & (new_n3992_ | new_n3449_ | new_n3444_ | ~P3_STATE2_REG_1__SCAN_IN);
  assign new_n3990_ = ~new_n3991_ & (~new_n3450_ ^ P3_PHYADDRPOINTER_REG_25__SCAN_IN) & (~P3_PHYADDRPOINTER_REG_30__SCAN_IN ^ (P3_PHYADDRPOINTER_REG_28__SCAN_IN & P3_PHYADDRPOINTER_REG_29__SCAN_IN & P3_PHYADDRPOINTER_REG_27__SCAN_IN & P3_PHYADDRPOINTER_REG_26__SCAN_IN & new_n3450_ & P3_PHYADDRPOINTER_REG_25__SCAN_IN));
  assign new_n3991_ = P3_PHYADDRPOINTER_REG_10__SCAN_IN ^ (new_n3334_ & P3_PHYADDRPOINTER_REG_9__SCAN_IN & P3_PHYADDRPOINTER_REG_7__SCAN_IN & P3_PHYADDRPOINTER_REG_8__SCAN_IN);
  assign new_n3992_ = (~new_n3334_ ^ P3_PHYADDRPOINTER_REG_7__SCAN_IN) & P3_PHYADDRPOINTER_REG_1__SCAN_IN & (~P3_PHYADDRPOINTER_REG_2__SCAN_IN ^ P3_PHYADDRPOINTER_REG_3__SCAN_IN);
  assign new_n3993_ = (~new_n2937_ | (~new_n3994_ & new_n3995_)) & (~P3_INSTADDRPOINTER_REG_1__SCAN_IN | new_n2937_ | new_n3282_) & (~P3_REIP_REG_1__SCAN_IN | P3_STATE2_REG_2__SCAN_IN | (~new_n2937_ & ~new_n3282_));
  assign new_n3994_ = (new_n2850_ | ~new_n3286_) & (~P3_INSTADDRPOINTER_REG_0__SCAN_IN | ~P3_INSTADDRPOINTER_REG_1__SCAN_IN) & (P3_INSTADDRPOINTER_REG_0__SCAN_IN | P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  assign new_n3995_ = (new_n3287_ | P3_INSTADDRPOINTER_REG_1__SCAN_IN) & (~new_n2928_ | new_n3927_) & (~new_n2927_ | new_n3928_);
  assign new_n3996_ = (new_n3471_ | new_n4005_) & ~new_n3998_ & (new_n4006_ | new_n3997_ | P3_STATE2_REG_2__SCAN_IN);
  assign new_n3997_ = ~new_n2937_ & ~new_n3282_;
  assign new_n3998_ = ((P3_EAX_REG_11__SCAN_IN & new_n3565_ & new_n3999_) | (new_n3565_ & ~new_n2826_) | (~P3_EAX_REG_11__SCAN_IN & (~new_n3565_ | ~new_n3999_))) & (new_n4000_ | ~new_n3565_ | ~new_n3522_) & (~BUF2_REG_11__SCAN_IN | new_n3522_ | ~new_n3565_ | new_n2826_);
  assign new_n3999_ = P3_EAX_REG_9__SCAN_IN & P3_EAX_REG_10__SCAN_IN & new_n3570_ & P3_EAX_REG_8__SCAN_IN;
  assign new_n4000_ = new_n4002_ & new_n4003_ & new_n4004_ & new_n4001_ & (~new_n2868_ | ~P3_INSTQUEUE_REG_0__3__SCAN_IN) & (~new_n2803_ | ~P3_INSTQUEUE_REG_9__3__SCAN_IN);
  assign new_n4001_ = (~P3_INSTQUEUE_REG_1__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P3_INSTQUEUE_REG_8__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_14__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n4002_ = (~P3_INSTQUEUE_REG_6__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_2__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_7__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n4003_ = (~P3_INSTQUEUE_REG_13__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_11__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_15__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_10__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n4004_ = (~P3_INSTQUEUE_REG_12__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P3_INSTQUEUE_REG_4__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_3__3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (~P3_INSTQUEUE_REG_5__3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  assign new_n4005_ = ~P3_EBX_REG_1__SCAN_IN & ~P3_EBX_REG_3__SCAN_IN & ~P3_EBX_REG_7__SCAN_IN & ~P3_EBX_REG_10__SCAN_IN & ~P3_EBX_REG_25__SCAN_IN & ~P3_EBX_REG_30__SCAN_IN;
  assign new_n4006_ = ~P3_REIP_REG_25__SCAN_IN & ~P3_REIP_REG_30__SCAN_IN & ~P3_REIP_REG_31__SCAN_IN & ~P3_REIP_REG_3__SCAN_IN & ~P3_REIP_REG_23__SCAN_IN;
  assign new_n4007_ = ~new_n4012_ & (new_n4014_ | ~new_n4015_) & new_n4008_ & (new_n2005_ | ~new_n2022_ | (~P2_REIP_REG_13__SCAN_IN & ~P2_REIP_REG_17__SCAN_IN));
  assign new_n4008_ = (~BUF2_REG_28__SCAN_IN | ~new_n3912_ | new_n2790_) & (~new_n4009_ | (new_n4011_ & new_n3915_)) & (~new_n4010_ | (new_n4011_ & P3_REIP_REG_1__SCAN_IN));
  assign new_n4009_ = new_n3910_ & new_n3472_ & P3_STATE2_REG_2__SCAN_IN & (~new_n3448_ | (new_n3445_ & ~new_n3447_));
  assign new_n4010_ = new_n3474_ & new_n3473_ & P3_STATE2_REG_2__SCAN_IN & (~new_n3448_ | (new_n3445_ & ~new_n3447_));
  assign new_n4011_ = P3_REIP_REG_30__SCAN_IN ^ (~P3_REIP_REG_28__SCAN_IN | ~P3_REIP_REG_29__SCAN_IN | ~new_n3484_ | ~P3_REIP_REG_27__SCAN_IN);
  assign new_n4012_ = ~new_n4013_ & (new_n2006_ | (~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_0__SCAN_IN & (~P2_STATE2_REG_2__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN))) & ((P2_STATE2_REG_2__SCAN_IN & ~P2_STATE2_REG_0__SCAN_IN) | (P2_STATE2_REG_1__SCAN_IN & ~P2_STATEBS16_REG_SCAN_IN));
  assign new_n4013_ = (~new_n2745_ ^ P2_PHYADDRPOINTER_REG_13__SCAN_IN) & (~new_n2018_ ^ P2_PHYADDRPOINTER_REG_17__SCAN_IN);
  assign new_n4014_ = (((P3_INSTADDRPOINTER_REG_4__SCAN_IN | (new_n2866_ ^ ~new_n2889_)) & (new_n2905_ | (P3_INSTADDRPOINTER_REG_4__SCAN_IN & (~new_n2866_ | new_n2889_) & (new_n2866_ | ~new_n2889_)))) | (P3_INSTADDRPOINTER_REG_5__SCAN_IN ^ (~new_n2894_ ^ (new_n2866_ & ~new_n2889_)))) & new_n3306_ & ((~P3_INSTADDRPOINTER_REG_4__SCAN_IN & (~new_n2866_ ^ ~new_n2889_)) | (~new_n2905_ & (~P3_INSTADDRPOINTER_REG_4__SCAN_IN | (new_n2866_ & ~new_n2889_) | (~new_n2866_ & new_n2889_))) | (P3_INSTADDRPOINTER_REG_5__SCAN_IN & (new_n2894_ | ~new_n2866_ | new_n2889_) & (~new_n2894_ | (new_n2866_ & ~new_n2889_))) | (~P3_INSTADDRPOINTER_REG_5__SCAN_IN & (new_n2894_ ^ (new_n2866_ & ~new_n2889_))));
  assign new_n4015_ = ~new_n4017_ & ~new_n4018_ & ~new_n4020_ & (new_n3296_ | ~new_n4022_) & ((new_n4016_ & new_n4021_) | ~new_n3332_ | (~new_n4016_ & ~new_n4021_));
  assign new_n4016_ = (new_n2918_ | ~new_n2920_) & (new_n2917_ | P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  assign new_n4017_ = P3_REIP_REG_5__SCAN_IN & new_n3284_ & (new_n3294_ | (new_n2950_ & ((new_n2927_ & new_n2939_) | (new_n2928_ & new_n2945_))));
  assign new_n4018_ = new_n4019_ & new_n3305_ & (new_n3294_ | (new_n2950_ & ((new_n2927_ & new_n2939_) | (new_n2928_ & new_n2945_))));
  assign new_n4019_ = P3_PHYADDRPOINTER_REG_5__SCAN_IN ^ (P3_PHYADDRPOINTER_REG_4__SCAN_IN & P3_PHYADDRPOINTER_REG_2__SCAN_IN & P3_PHYADDRPOINTER_REG_3__SCAN_IN);
  assign new_n4020_ = P3_PHYADDRPOINTER_REG_5__SCAN_IN & ~new_n3294_ & (~new_n2950_ | ((~new_n2927_ | ~new_n2939_) & (~new_n2928_ | ~new_n2945_)));
  assign new_n4021_ = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN ^ (new_n2894_ ^ (~new_n2889_ & ~new_n2878_ & ~new_n2867_ & ~new_n2873_));
  assign new_n4022_ = (~P3_PHYADDRPOINTER_REG_1__SCAN_IN | ~P3_PHYADDRPOINTER_REG_5__SCAN_IN | ~P3_PHYADDRPOINTER_REG_4__SCAN_IN | ~P3_PHYADDRPOINTER_REG_2__SCAN_IN | ~P3_PHYADDRPOINTER_REG_3__SCAN_IN) & (P3_PHYADDRPOINTER_REG_5__SCAN_IN | (P3_PHYADDRPOINTER_REG_1__SCAN_IN & P3_PHYADDRPOINTER_REG_4__SCAN_IN & P3_PHYADDRPOINTER_REG_2__SCAN_IN & P3_PHYADDRPOINTER_REG_3__SCAN_IN));
  assign new_n4023_ = new_n3443_ & (~P3_PHYADDRPOINTER_REG_10__SCAN_IN | ~new_n3334_ | ~P3_PHYADDRPOINTER_REG_9__SCAN_IN | ~P3_PHYADDRPOINTER_REG_7__SCAN_IN | ~P3_PHYADDRPOINTER_REG_8__SCAN_IN | P3_PHYADDRPOINTER_REG_0__SCAN_IN | ~P3_PHYADDRPOINTER_REG_1__SCAN_IN) & ((P3_PHYADDRPOINTER_REG_10__SCAN_IN & new_n3334_ & P3_PHYADDRPOINTER_REG_9__SCAN_IN & P3_PHYADDRPOINTER_REG_7__SCAN_IN & P3_PHYADDRPOINTER_REG_8__SCAN_IN) | (~P3_PHYADDRPOINTER_REG_10__SCAN_IN & (~new_n3334_ | ~P3_PHYADDRPOINTER_REG_9__SCAN_IN | ~P3_PHYADDRPOINTER_REG_7__SCAN_IN | ~P3_PHYADDRPOINTER_REG_8__SCAN_IN)) | (~P3_PHYADDRPOINTER_REG_10__SCAN_IN & ~P3_PHYADDRPOINTER_REG_0__SCAN_IN & P3_PHYADDRPOINTER_REG_1__SCAN_IN & P3_PHYADDRPOINTER_REG_8__SCAN_IN & new_n3334_ & P3_PHYADDRPOINTER_REG_7__SCAN_IN));
  assign new_n4024_ = new_n4025_ & new_n4028_ & new_n4039_ & ~new_n2636_ & ~new_n4030_ & new_n4032_;
  assign new_n4025_ = (~new_n4026_ | ~new_n2585_ | ~new_n2495_ | (~new_n2566_ & new_n2568_)) & (~new_n4027_ | new_n2572_ | ~new_n2495_ | (~new_n2566_ & new_n2568_));
  assign new_n4026_ = P1_INSTADDRPOINTER_REG_20__SCAN_IN ^ (new_n2583_ & P1_INSTADDRPOINTER_REG_17__SCAN_IN & P1_INSTADDRPOINTER_REG_16__SCAN_IN & P1_INSTADDRPOINTER_REG_15__SCAN_IN & new_n2579_ & P1_INSTADDRPOINTER_REG_14__SCAN_IN);
  assign new_n4027_ = new_n2470_ ^ (new_n2454_ & ~new_n2469_ & new_n2468_ & new_n2467_ & new_n2457_ & new_n2463_);
  assign new_n4028_ = (~new_n2585_ | ~new_n2495_ | (~new_n2566_ & new_n2568_) | (new_n2579_ & P1_INSTADDRPOINTER_REG_14__SCAN_IN) | (~new_n2579_ & ~P1_INSTADDRPOINTER_REG_14__SCAN_IN)) & (new_n4029_ | ~new_n2493_ | ~new_n2495_ | (~new_n2566_ & new_n2568_));
  assign new_n4029_ = (~new_n2592_ ^ P1_INSTADDRPOINTER_REG_17__SCAN_IN) & (~P1_INSTADDRPOINTER_REG_20__SCAN_IN ^ (new_n2583_ & new_n2592_ & P1_INSTADDRPOINTER_REG_17__SCAN_IN));
  assign new_n4030_ = ~P2_STATE2_REG_2__SCAN_IN & (new_n2706_ | new_n4031_) & (P2_REIP_REG_7__SCAN_IN | P2_REIP_REG_2__SCAN_IN | P2_REIP_REG_5__SCAN_IN);
  assign new_n4031_ = new_n2022_ & ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_0__SCAN_IN;
  assign new_n4032_ = (~new_n3502_ | (~P1_REIP_REG_21__SCAN_IN & ~P1_REIP_REG_6__SCAN_IN)) & (new_n4033_ | new_n4035_ | ~new_n4036_ | (~new_n3471_ & P3_EBX_REG_8__SCAN_IN));
  assign new_n4033_ = new_n3449_ & ~new_n3444_ & P3_STATE2_REG_1__SCAN_IN & (P3_PHYADDRPOINTER_REG_0__SCAN_IN | ~P3_PHYADDRPOINTER_REG_1__SCAN_IN | ~new_n4034_ | ~P3_PHYADDRPOINTER_REG_8__SCAN_IN) & ((new_n4034_ & P3_PHYADDRPOINTER_REG_8__SCAN_IN) | (~new_n4034_ & ~P3_PHYADDRPOINTER_REG_8__SCAN_IN) | (new_n4034_ & ~P3_PHYADDRPOINTER_REG_0__SCAN_IN & P3_PHYADDRPOINTER_REG_1__SCAN_IN));
  assign new_n4034_ = new_n3334_ & P3_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign new_n4035_ = ~new_n3449_ & ~new_n3444_ & P3_STATE2_REG_1__SCAN_IN & (new_n4034_ | P3_PHYADDRPOINTER_REG_8__SCAN_IN) & (~new_n4034_ | ~P3_PHYADDRPOINTER_REG_8__SCAN_IN);
  assign new_n4036_ = (~new_n3476_ | (~new_n3480_ & P3_EBX_REG_8__SCAN_IN) | (new_n3480_ & ~P3_EBX_REG_8__SCAN_IN)) & (new_n3483_ | ~new_n4038_) & new_n4037_ & (~new_n3498_ | ~P3_PHYADDRPOINTER_REG_8__SCAN_IN);
  assign new_n4037_ = (new_n3448_ & (~new_n3445_ | new_n3447_)) ? ~P3_REIP_REG_8__SCAN_IN : (P3_STATE2_REG_1__SCAN_IN | P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN);
  assign new_n4038_ = ~P3_REIP_REG_8__SCAN_IN ^ (~new_n3916_ | ~P3_REIP_REG_7__SCAN_IN);
  assign new_n4039_ = ~new_n4040_ & (~new_n2509_ | ((~new_n3349_ | ~new_n2067_ | (~P1_EAX_REG_11__SCAN_IN & ~P1_EAX_REG_8__SCAN_IN)) & (~new_n4041_ | ~new_n3349_ | new_n2067_)));
  assign new_n4040_ = (P3_INSTADDRPOINTER_REG_21__SCAN_IN | (P3_INSTADDRPOINTER_REG_20__SCAN_IN & P3_INSTADDRPOINTER_REG_19__SCAN_IN & new_n2781_ & new_n2924_ & (new_n2913_ | ~new_n2922_))) & new_n3307_ & (~P3_INSTADDRPOINTER_REG_21__SCAN_IN | ~P3_INSTADDRPOINTER_REG_20__SCAN_IN | ~P3_INSTADDRPOINTER_REG_19__SCAN_IN | ~new_n2781_ | ~new_n2924_ | (~new_n2913_ & new_n2922_));
  assign new_n4041_ = new_n2954_ ? (BUF1_REG_8__SCAN_IN | BUF1_REG_11__SCAN_IN) : (DATAI_11_ | DATAI_8_);
  assign new_n4042_ = new_n4051_ & new_n4066_ & new_n4043_ & new_n4049_;
  assign new_n4043_ = (~new_n2589_ | ~P1_REIP_REG_14__SCAN_IN) & ~new_n4044_ & ~new_n4048_ & ((P3_INSTADDRPOINTER_REG_16__SCAN_IN & new_n3291_ & P3_INSTADDRPOINTER_REG_15__SCAN_IN) | ~new_n3307_ | (~P3_INSTADDRPOINTER_REG_16__SCAN_IN & (~new_n3291_ | ~P3_INSTADDRPOINTER_REG_15__SCAN_IN)));
  assign new_n4044_ = (~new_n4045_ | P2_STATE2_REG_0__SCAN_IN | (~new_n3439_ & (~P2_STATE2_REG_2__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN))) & (~new_n4046_ | new_n3439_ | (P2_STATE2_REG_1__SCAN_IN & P2_STATE2_REG_2__SCAN_IN & ~P2_STATE2_REG_0__SCAN_IN)) & (~new_n3439_ | ~new_n4047_ | ~P2_STATE2_REG_0__SCAN_IN | ~P2_EAX_REG_3__SCAN_IN);
  assign new_n4045_ = P2_LWORD_REG_3__SCAN_IN & P2_LWORD_REG_14__SCAN_IN & P2_LWORD_REG_8__SCAN_IN;
  assign new_n4046_ = P2_DATAO_REG_14__SCAN_IN & P2_DATAO_REG_3__SCAN_IN & P2_DATAO_REG_8__SCAN_IN;
  assign new_n4047_ = P2_EAX_REG_8__SCAN_IN & P2_EAX_REG_14__SCAN_IN;
  assign new_n4048_ = (~P1_UWORD_REG_0__SCAN_IN | P1_STATE2_REG_0__SCAN_IN | (~new_n3509_ & ~new_n3312_)) & (~P1_EAX_REG_16__SCAN_IN | ~new_n3509_ | new_n2073_ | ~P1_STATE2_REG_0__SCAN_IN) & (~P1_DATAO_REG_16__SCAN_IN | new_n3509_ | new_n3312_);
  assign new_n4049_ = ~new_n4050_ & (new_n2630_ | ~P1_STATE2_REG_3__SCAN_IN | (~P1_PHYADDRPOINTER_REG_23__SCAN_IN & ~P1_PHYADDRPOINTER_REG_22__SCAN_IN & ~P1_PHYADDRPOINTER_REG_4__SCAN_IN & ~P1_PHYADDRPOINTER_REG_19__SCAN_IN & ~P1_PHYADDRPOINTER_REG_12__SCAN_IN));
  assign new_n4050_ = (~P1_LWORD_REG_3__SCAN_IN | (new_n3349_ & new_n2509_)) & (~new_n2509_ | ((~P1_EAX_REG_3__SCAN_IN | ~new_n3349_ | ~new_n2067_) & (~new_n3349_ | new_n2067_ | (new_n2954_ ? ~BUF1_REG_3__SCAN_IN : ~DATAI_3_))));
  assign new_n4051_ = new_n4052_ & new_n4053_ & ~new_n4064_ & ~new_n4065_ & new_n4054_ & new_n4060_ & new_n4061_;
  assign new_n4052_ = (~new_n3095_ | new_n2091_ | ~P1_STATE2_REG_3__SCAN_IN | P1_STATE2_REG_0__SCAN_IN | (~new_n2997_ & (new_n2477_ | ~P1_STATE2_REG_3__SCAN_IN))) & (~new_n3042_ | new_n2067_ | ~P1_STATE2_REG_3__SCAN_IN | P1_STATE2_REG_0__SCAN_IN | (~new_n2997_ & (new_n2477_ | ~P1_STATE2_REG_3__SCAN_IN)));
  assign new_n4053_ = (~new_n3017_ | new_n2079_ | ~P1_STATE2_REG_3__SCAN_IN | P1_STATE2_REG_0__SCAN_IN | (~new_n2997_ & (new_n2477_ | ~P1_STATE2_REG_3__SCAN_IN))) & (~new_n3219_ | new_n2065_ | ~P1_STATE2_REG_3__SCAN_IN | P1_STATE2_REG_0__SCAN_IN | (~new_n2997_ & (new_n2477_ | ~P1_STATE2_REG_3__SCAN_IN)));
  assign new_n4054_ = (~new_n4056_ | ~new_n2706_ | new_n4055_) & ((new_n4056_ & ~new_n4057_) | ~new_n2706_ | ~new_n1783_) & (new_n4058_ | new_n2706_ | new_n4031_) & (~new_n4059_ | ~new_n2706_ | new_n4055_);
  assign new_n4055_ = new_n3172_ & (~new_n1760_ | new_n1322_ | new_n1370_) & (~new_n2708_ | new_n1322_ | ~new_n1370_);
  assign new_n4056_ = ~P2_INSTADDRPOINTER_REG_2__SCAN_IN ^ (~P2_INSTADDRPOINTER_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_1__SCAN_IN);
  assign new_n4057_ = P2_INSTADDRPOINTER_REG_5__SCAN_IN ^ (P2_INSTADDRPOINTER_REG_3__SCAN_IN & P2_INSTADDRPOINTER_REG_4__SCAN_IN & (P2_INSTADDRPOINTER_REG_2__SCAN_IN | (P2_INSTADDRPOINTER_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_1__SCAN_IN)));
  assign new_n4058_ = ~P2_INSTADDRPOINTER_REG_7__SCAN_IN & ~P2_INSTADDRPOINTER_REG_2__SCAN_IN & ~P2_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign new_n4059_ = (~P2_INSTADDRPOINTER_REG_7__SCAN_IN | ~P2_INSTADDRPOINTER_REG_6__SCAN_IN | ~P2_INSTADDRPOINTER_REG_5__SCAN_IN | ~P2_INSTADDRPOINTER_REG_3__SCAN_IN | ~P2_INSTADDRPOINTER_REG_4__SCAN_IN | ~P2_INSTADDRPOINTER_REG_2__SCAN_IN | ~P2_INSTADDRPOINTER_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_1__SCAN_IN) & ((P2_INSTADDRPOINTER_REG_5__SCAN_IN ^ (P2_INSTADDRPOINTER_REG_3__SCAN_IN & P2_INSTADDRPOINTER_REG_4__SCAN_IN & P2_INSTADDRPOINTER_REG_2__SCAN_IN & P2_INSTADDRPOINTER_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_1__SCAN_IN)) | P2_INSTADDRPOINTER_REG_7__SCAN_IN | (P2_INSTADDRPOINTER_REG_6__SCAN_IN & P2_INSTADDRPOINTER_REG_5__SCAN_IN & P2_INSTADDRPOINTER_REG_3__SCAN_IN & P2_INSTADDRPOINTER_REG_4__SCAN_IN & P2_INSTADDRPOINTER_REG_2__SCAN_IN & P2_INSTADDRPOINTER_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_1__SCAN_IN));
  assign new_n4060_ = (new_n1335_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (new_n1367_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  assign new_n4061_ = (~new_n2706_ | new_n4062_ | (new_n1387_ & ~new_n1410_) | (~new_n1387_ & new_n1410_)) & (~new_n2706_ | ~new_n1783_ | (~new_n4063_ & ~P2_INSTADDRPOINTER_REG_7__SCAN_IN) | (new_n4063_ & P2_INSTADDRPOINTER_REG_7__SCAN_IN));
  assign new_n4062_ = (~new_n1322_ | new_n1335_ | new_n1317_ | new_n1330_ | ~new_n1350_ | ~new_n1370_ | ~new_n1345_ | new_n1367_) & (~new_n1322_ | new_n1370_ | ~new_n1350_ | new_n1335_ | new_n1345_ | ~new_n1330_ | ~new_n1317_ | ~new_n1367_) & (~new_n1345_ | ~new_n1367_ | ~new_n1330_ | new_n1335_ | ~new_n1322_ | new_n1317_ | ~new_n1370_) & (~new_n1345_ | ~new_n1367_ | ~new_n1330_ | new_n1335_ | new_n1350_ | ~new_n1317_ | ~new_n1322_ | ~new_n1370_);
  assign new_n4063_ = P2_INSTADDRPOINTER_REG_6__SCAN_IN & P2_INSTADDRPOINTER_REG_5__SCAN_IN & P2_INSTADDRPOINTER_REG_3__SCAN_IN & P2_INSTADDRPOINTER_REG_4__SCAN_IN & (P2_INSTADDRPOINTER_REG_2__SCAN_IN | (P2_INSTADDRPOINTER_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_1__SCAN_IN));
  assign new_n4064_ = (~new_n3509_ | ~P1_EAX_REG_10__SCAN_IN) & (~P1_DATAO_REG_10__SCAN_IN | new_n3509_ | new_n3312_) & (~P1_LWORD_REG_10__SCAN_IN | P1_STATE2_REG_0__SCAN_IN | (~new_n3509_ & ~new_n3312_));
  assign new_n4065_ = new_n3013_ & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n4066_ = new_n4067_ & (~new_n3013_ | ~new_n3223_) & (new_n2505_ | ~P1_EAX_REG_16__SCAN_IN) & new_n4069_ & ~new_n4070_ & (new_n2505_ | ~P1_EAX_REG_23__SCAN_IN);
  assign new_n4067_ = (~new_n4068_ | ~new_n3037_) & ((P1_LWORD_REG_1__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN & (new_n3509_ | new_n3312_)) | (new_n3509_ & P1_EAX_REG_1__SCAN_IN) | (P1_DATAO_REG_1__SCAN_IN & ~new_n3509_ & ~new_n3312_));
  assign new_n4068_ = ~new_n2053_ & P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN & (new_n2997_ | (P1_STATE2_REG_3__SCAN_IN & (new_n2478_ | new_n2482_)));
  assign new_n4069_ = (~new_n4068_ | ((P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN))) & (~new_n3351_ | P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  assign new_n4070_ = new_n3351_ & new_n3095_;
  assign new_n4071_ = ~new_n4072_ & ~new_n4075_ & ~new_n4079_ & (~new_n4078_ | (~new_n3313_ & (~new_n1978_ ^ ~new_n1984_)));
  assign new_n4072_ = new_n2756_ & (~new_n4073_ | (new_n2728_ ^ P2_PHYADDRPOINTER_REG_31__SCAN_IN));
  assign new_n4073_ = (~new_n2016_ ^ P2_PHYADDRPOINTER_REG_25__SCAN_IN) & new_n4074_ & (P2_PHYADDRPOINTER_REG_22__SCAN_IN ^ (~new_n2731_ | ~P2_PHYADDRPOINTER_REG_21__SCAN_IN));
  assign new_n4074_ = (~P2_PHYADDRPOINTER_REG_20__SCAN_IN ^ (P2_PHYADDRPOINTER_REG_19__SCAN_IN & new_n2732_ & P2_PHYADDRPOINTER_REG_18__SCAN_IN)) & (new_n2745_ ^ ~P2_PHYADDRPOINTER_REG_13__SCAN_IN) & (~P2_PHYADDRPOINTER_REG_15__SCAN_IN ^ (P2_PHYADDRPOINTER_REG_14__SCAN_IN & new_n2745_ & P2_PHYADDRPOINTER_REG_13__SCAN_IN));
  assign new_n4075_ = ~new_n4076_ & P1_EBX_REG_31__SCAN_IN & ~new_n2634_ & ~new_n2630_ & new_n2494_ & P1_STATE2_REG_2__SCAN_IN;
  assign new_n4076_ = (~new_n2453_ ^ new_n2473_) & (~new_n2467_ ^ (new_n2457_ & new_n2463_)) & ~new_n3262_ & (new_n2770_ ^ new_n4077_);
  assign new_n4077_ = new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_4__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_4__SCAN_IN));
  assign new_n4078_ = new_n2706_ & ~new_n4062_;
  assign new_n4079_ = (~P3_INSTADDRPOINTER_REG_16__SCAN_IN | ~P3_INSTADDRPOINTER_REG_15__SCAN_IN | ~new_n3278_ | ~new_n2782_) & new_n3306_ & (P3_INSTADDRPOINTER_REG_16__SCAN_IN | (P3_INSTADDRPOINTER_REG_15__SCAN_IN & new_n3278_ & new_n2782_));
  assign new_n4080_ = new_n4087_ & new_n4088_ & new_n4081_ & new_n4082_;
  assign new_n4081_ = (~new_n3188_ | ~new_n2963_ | (new_n1664_ & (~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_))) | (~new_n1664_ & ((new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_)))) | (~new_n1412_ & (new_n1409_ | ~new_n1421_) & (~new_n1409_ | new_n1421_)) | (new_n1412_ & (new_n1409_ ^ new_n1421_))) & (~new_n3069_ | ~new_n3059_ | (new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) | (~new_n1412_ ^ (~new_n1409_ ^ new_n1421_)));
  assign new_n4082_ = ~new_n4084_ & (~new_n4083_ | ~new_n2963_ | (new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) | (~new_n1412_ & (~new_n1409_ | new_n1421_) & (new_n1409_ | ~new_n1421_)) | (new_n1412_ & (~new_n1409_ ^ ~new_n1421_)));
  assign new_n4083_ = new_n2968_ & (new_n2976_ ? BUF1_REG_31__SCAN_IN : BUF2_REG_31__SCAN_IN);
  assign new_n4084_ = ~new_n4085_ & new_n2644_ & new_n2275_ & P1_STATE2_REG_1__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN;
  assign new_n4085_ = (~P1_PHYADDRPOINTER_REG_23__SCAN_IN ^ (P1_PHYADDRPOINTER_REG_22__SCAN_IN & P1_PHYADDRPOINTER_REG_21__SCAN_IN & new_n2354_ & P1_PHYADDRPOINTER_REG_20__SCAN_IN)) & new_n4086_ & (~P1_PHYADDRPOINTER_REG_22__SCAN_IN ^ (P1_PHYADDRPOINTER_REG_21__SCAN_IN & new_n2354_ & P1_PHYADDRPOINTER_REG_20__SCAN_IN));
  assign new_n4086_ = ~new_n2366_ & ~new_n2246_ & P1_PHYADDRPOINTER_REG_1__SCAN_IN & (~P1_PHYADDRPOINTER_REG_4__SCAN_IN ^ (P1_PHYADDRPOINTER_REG_3__SCAN_IN & P1_PHYADDRPOINTER_REG_2__SCAN_IN & P1_PHYADDRPOINTER_REG_1__SCAN_IN));
  assign new_n4087_ = (~new_n3244_ | ~new_n2963_ | (new_n1664_ & (~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_))) | (~new_n1664_ & ((new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_)))) | (~new_n1412_ & (new_n1409_ | ~new_n1421_) & (~new_n1409_ | new_n1421_)) | (new_n1412_ & (new_n1409_ ^ new_n1421_))) & (~new_n3241_ | new_n1666_ | (new_n1664_ & (~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_))) | (~new_n1664_ & ((new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_)))) | (~new_n1412_ & (new_n1409_ | ~new_n1421_) & (~new_n1409_ | new_n1421_)) | (new_n1412_ & (new_n1409_ ^ new_n1421_)));
  assign new_n4088_ = (~new_n2968_ | new_n3194_ | ~new_n2963_ | (new_n1664_ & (~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_))) | (~new_n1664_ & ((new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_)))) | (~new_n1412_ ^ (~new_n1409_ ^ new_n1421_))) & (~new_n2968_ | ~new_n3210_ | ~new_n2963_ | (new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) | (~new_n1412_ ^ (~new_n1409_ ^ new_n1421_)));
  assign new_n4089_ = new_n4097_ & (~new_n4095_ | (new_n2726_ & new_n4099_) | ~new_n4090_ | (~new_n2723_ & P2_EBX_REG_4__SCAN_IN));
  assign new_n4090_ = ((new_n1981_ & (new_n4093_ | new_n4094_) & (new_n4092_ | (new_n4093_ & new_n4094_))) | ~new_n2691_ | (~new_n1981_ & ((~new_n4093_ & ~new_n4094_) | (~new_n4092_ & (~new_n4093_ | ~new_n4094_))))) & new_n4091_ & (~new_n1891_ | ~new_n2757_);
  assign new_n4091_ = (~new_n2665_ | ~new_n1673_) & (~P2_PHYADDRPOINTER_REG_4__SCAN_IN | new_n2724_ | ~P2_STATE2_REG_3__SCAN_IN) & (~new_n2724_ | ~P2_REIP_REG_4__SCAN_IN) & (new_n2724_ | ~new_n3374_);
  assign new_n4092_ = ~new_n1383_ & (new_n1386_ | new_n1387_);
  assign new_n4093_ = (~new_n1382_ | ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | (new_n1328_ & new_n1365_));
  assign new_n4094_ = new_n1379_ & (new_n1373_ | ~P2_INSTADDRPOINTER_REG_3__SCAN_IN);
  assign new_n4095_ = (~new_n4096_ | (new_n1662_ & new_n1420_) | (~new_n1662_ & ~new_n1420_)) & (~new_n2756_ | (P2_PHYADDRPOINTER_REG_4__SCAN_IN & P2_PHYADDRPOINTER_REG_3__SCAN_IN & P2_PHYADDRPOINTER_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_2__SCAN_IN) | (~P2_PHYADDRPOINTER_REG_4__SCAN_IN & (~P2_PHYADDRPOINTER_REG_3__SCAN_IN | ~P2_PHYADDRPOINTER_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_2__SCAN_IN)));
  assign new_n4096_ = new_n1370_ & new_n2666_ & P2_STATE2_REG_2__SCAN_IN;
  assign new_n4097_ = (~new_n4098_ | ~new_n3012_) & (~new_n4098_ | new_n3270_);
  assign new_n4098_ = (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & new_n2284_ & new_n2994_ & (new_n2154_ | (new_n2148_ & new_n2200_) | (~new_n2148_ & ~new_n2200_)) & (~new_n2154_ | (new_n2148_ ^ new_n2200_));
  assign new_n4099_ = (P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_4__SCAN_IN : (~P2_PHYADDRPOINTER_REG_4__SCAN_IN ^ (P2_PHYADDRPOINTER_REG_3__SCAN_IN & P2_PHYADDRPOINTER_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_2__SCAN_IN))) ^ (new_n2740_ & (~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_3__SCAN_IN) & ((~P2_PHYADDRPOINTER_REG_3__SCAN_IN & (~P2_PHYADDRPOINTER_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_2__SCAN_IN)) | P2_STATE2_REG_0__SCAN_IN | (P2_PHYADDRPOINTER_REG_3__SCAN_IN & P2_PHYADDRPOINTER_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_2__SCAN_IN)));
  assign new_n4100_ = ~new_n4117_ & ((P3_STATE2_REG_1__SCAN_IN & (((new_n4101_ | ~P3_STATE2_REG_0__SCAN_IN) & P3_STATE2_REG_2__SCAN_IN & (P3_STATE2_REG_0__SCAN_IN | (new_n2943_ & P3_STATE2_REG_1__SCAN_IN))) | (new_n2943_ & ~P3_STATE2_REG_2__SCAN_IN & P3_STATE2_REG_0__SCAN_IN))) | (((~new_n4101_ & P3_STATE2_REG_0__SCAN_IN) | ~P3_STATE2_REG_2__SCAN_IN | (~P3_STATE2_REG_0__SCAN_IN & (~new_n2943_ | ~P3_STATE2_REG_1__SCAN_IN))) & ((P3_STATE2_REG_0__SCAN_IN & P3_STATE2_REG_2__SCAN_IN & ~P3_STATE2_REG_1__SCAN_IN) | (~P3_STATE2_REG_3__SCAN_IN & ~P3_STATE2_REG_1__SCAN_IN & ~new_n2943_ & P3_STATE2_REG_0__SCAN_IN))) | (~P3_STATE2_REG_2__SCAN_IN & ~P3_STATE2_REG_0__SCAN_IN & P3_STATE2_REG_1__SCAN_IN & ~P3_STATEBS16_REG_SCAN_IN));
  assign new_n4101_ = (new_n4102_ | (new_n4113_ & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) | (~new_n4110_ & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN)) & (new_n4106_ | ~new_n4110_) & new_n4113_ & new_n4114_;
  assign new_n4102_ = ((~new_n4105_ & (new_n4103_ | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)) | (new_n4106_ & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) | (new_n4103_ & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)) & (new_n4106_ | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & (~new_n4110_ | P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  assign new_n4103_ = ((new_n3528_ & ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~new_n3525_ & new_n3526_) | new_n4104_ | (new_n3287_ & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN)) & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & (~new_n4104_ | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  assign new_n4104_ = ~new_n3517_ & new_n3519_ & new_n3521_;
  assign new_n4105_ = new_n4104_ ? P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN : ~new_n3524_;
  assign new_n4106_ = (new_n4104_ | new_n4107_) & (~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | (~new_n4104_ & ((new_n2861_ & new_n4109_) | (P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN))));
  assign new_n4107_ = ((~new_n4108_ & new_n3527_) | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (new_n3527_ | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~new_n2850_ | (P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ (P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN))) & (~new_n2832_ | (P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN));
  assign new_n4108_ = P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & (new_n2789_ | ~new_n3526_);
  assign new_n4109_ = (~new_n2826_ | ~new_n2821_ | ~new_n2833_ | new_n2790_ | new_n2796_ | new_n2815_ | new_n2802_ | ~new_n2809_) & (new_n2802_ | ~new_n2833_ | new_n2790_ | new_n2796_ | ~new_n2815_ | new_n2826_ | new_n2821_) & ((new_n2802_ ^ new_n2809_) | ~new_n2826_ | ~new_n2833_ | ~new_n2815_ | ~new_n2821_ | new_n2790_ | ~new_n2796_) & (~new_n2802_ | ~new_n2790_ | ~new_n2821_ | ((~new_n2815_ | new_n2833_) & (~new_n2826_ | ~new_n2833_ | ~new_n2796_ | new_n2815_)));
  assign new_n4110_ = (~new_n4104_ | P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~new_n4111_ | ((P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | (new_n3922_ & (new_n4108_ | ~new_n3287_))) & (new_n4104_ | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | (~new_n4112_ & (~new_n2861_ | (~new_n3287_ & ~new_n3922_))))));
  assign new_n4111_ = (new_n4109_ | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | (P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN)) & (~new_n2850_ | (P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN & (P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | (P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN))) | (~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN & (~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN)));
  assign new_n4112_ = P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign new_n4113_ = new_n4104_ ? ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN : (~new_n2832_ | (new_n3921_ & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN) | (~new_n3921_ & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN));
  assign new_n4114_ = (new_n3581_ | new_n3824_) & (~new_n3581_ | (~P3_FLUSH_REG_SCAN_IN & ~P3_MORE_REG_SCAN_IN)) & ~new_n4115_ & ~P3_STATE2_REG_1__SCAN_IN & (~new_n3910_ | ~new_n3518_);
  assign new_n4115_ = (~new_n2802_ | new_n2945_) & new_n4116_ & ~new_n2809_ & (new_n2939_ | new_n2802_);
  assign new_n4116_ = new_n2833_ & ~new_n2790_ & ~new_n2796_ & new_n2815_ & ~new_n2826_ & ~new_n2821_;
  assign new_n4117_ = (~new_n2923_ | new_n2906_ | (~P3_INSTADDRPOINTER_REG_16__SCAN_IN ^ ((~P3_INSTADDRPOINTER_REG_15__SCAN_IN | (new_n2923_ & ~new_n2906_)) & ((~P3_INSTADDRPOINTER_REG_15__SCAN_IN & new_n2923_ & ~new_n2906_) | ((~P3_INSTADDRPOINTER_REG_14__SCAN_IN | (new_n2923_ & ~new_n2906_)) & (new_n2931_ | (~P3_INSTADDRPOINTER_REG_14__SCAN_IN & new_n2923_ & ~new_n2906_))))))) & new_n3332_ & ~new_n2906_ & (new_n2923_ | (~P3_INSTADDRPOINTER_REG_16__SCAN_IN & (~P3_INSTADDRPOINTER_REG_15__SCAN_IN | (new_n2923_ & ~new_n2906_)) & ((~P3_INSTADDRPOINTER_REG_15__SCAN_IN & new_n2923_ & ~new_n2906_) | ((~P3_INSTADDRPOINTER_REG_14__SCAN_IN | (new_n2923_ & ~new_n2906_)) & (new_n2931_ | (~P3_INSTADDRPOINTER_REG_14__SCAN_IN & new_n2923_ & ~new_n2906_))))) | (P3_INSTADDRPOINTER_REG_16__SCAN_IN & ((P3_INSTADDRPOINTER_REG_15__SCAN_IN & (~new_n2923_ | new_n2906_)) | ((P3_INSTADDRPOINTER_REG_15__SCAN_IN | ~new_n2923_ | new_n2906_) & ((P3_INSTADDRPOINTER_REG_14__SCAN_IN & (~new_n2923_ | new_n2906_)) | (~new_n2931_ & (P3_INSTADDRPOINTER_REG_14__SCAN_IN | ~new_n2923_ | new_n2906_)))))));
  assign new_n4118_ = ~new_n4119_ & (new_n4126_ | ~new_n4124_ | new_n4127_ | (new_n2756_ & (P2_PHYADDRPOINTER_REG_1__SCAN_IN | P2_PHYADDRPOINTER_REG_2__SCAN_IN) & (~P2_PHYADDRPOINTER_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_2__SCAN_IN)));
  assign new_n4119_ = ~new_n4120_ & ~new_n4121_ & ~new_n4122_ & (~new_n2665_ | ~new_n1676_) & new_n4123_ & (new_n2723_ | ~P2_EBX_REG_6__SCAN_IN);
  assign new_n4120_ = new_n2726_ & ((P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_6__SCAN_IN) | (~P2_STATE2_REG_0__SCAN_IN & (~P2_PHYADDRPOINTER_REG_6__SCAN_IN | ~new_n2743_ | ~P2_PHYADDRPOINTER_REG_5__SCAN_IN) & (P2_PHYADDRPOINTER_REG_6__SCAN_IN | (new_n2743_ & P2_PHYADDRPOINTER_REG_5__SCAN_IN))) | ~new_n2739_ | (P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_5__SCAN_IN) | (~P2_STATE2_REG_0__SCAN_IN & (~new_n2743_ | ~P2_PHYADDRPOINTER_REG_5__SCAN_IN) & (new_n2743_ | P2_PHYADDRPOINTER_REG_5__SCAN_IN))) & ((P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_6__SCAN_IN : (~P2_PHYADDRPOINTER_REG_6__SCAN_IN ^ (new_n2743_ & P2_PHYADDRPOINTER_REG_5__SCAN_IN))) | (new_n2739_ & (~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_5__SCAN_IN) & (P2_STATE2_REG_0__SCAN_IN | (new_n2743_ & P2_PHYADDRPOINTER_REG_5__SCAN_IN) | (~new_n2743_ & ~P2_PHYADDRPOINTER_REG_5__SCAN_IN))));
  assign new_n4121_ = new_n2756_ & (~P2_PHYADDRPOINTER_REG_6__SCAN_IN | ~new_n2743_ | ~P2_PHYADDRPOINTER_REG_5__SCAN_IN) & (P2_PHYADDRPOINTER_REG_6__SCAN_IN | (new_n2743_ & P2_PHYADDRPOINTER_REG_5__SCAN_IN));
  assign new_n4122_ = (~new_n1983_ | (~new_n1982_ & ~new_n1981_ & ((~new_n4093_ & ~new_n4094_) | (~new_n4092_ & (~new_n4093_ | ~new_n4094_))))) & new_n2691_ & (new_n1983_ | new_n1982_ | new_n1981_ | ((new_n4093_ | new_n4094_) & (new_n4092_ | (new_n4093_ & new_n4094_))));
  assign new_n4123_ = (~new_n2757_ | ~new_n1883_) & (~P2_PHYADDRPOINTER_REG_6__SCAN_IN | new_n2724_ | ~P2_STATE2_REG_3__SCAN_IN) & (~new_n2724_ | ~P2_REIP_REG_6__SCAN_IN) & (new_n2724_ | ~new_n3374_);
  assign new_n4124_ = (new_n2723_ | ~P2_EBX_REG_2__SCAN_IN) & new_n4125_ & (~new_n2757_ | ~new_n1902_);
  assign new_n4125_ = (~new_n1814_ | ~new_n2691_) & (~new_n2665_ | ~new_n1667_) & (~new_n2724_ | ~P2_REIP_REG_2__SCAN_IN) & (~P2_PHYADDRPOINTER_REG_2__SCAN_IN | new_n2724_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n4126_ = new_n2726_ & ((P2_STATE2_REG_0__SCAN_IN ? P2_INSTADDRPOINTER_REG_0__SCAN_IN : P2_PHYADDRPOINTER_REG_0__SCAN_IN) | (P2_STATE2_REG_0__SCAN_IN ? P2_INSTADDRPOINTER_REG_1__SCAN_IN : ~P2_PHYADDRPOINTER_REG_1__SCAN_IN) | (P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_2__SCAN_IN) | (~P2_STATE2_REG_0__SCAN_IN & (~P2_PHYADDRPOINTER_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_2__SCAN_IN) & (P2_PHYADDRPOINTER_REG_1__SCAN_IN | P2_PHYADDRPOINTER_REG_2__SCAN_IN))) & (((P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_0__SCAN_IN : ~P2_PHYADDRPOINTER_REG_0__SCAN_IN) & (P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_1__SCAN_IN : P2_PHYADDRPOINTER_REG_1__SCAN_IN)) | (P2_STATE2_REG_0__SCAN_IN ? ~P2_INSTADDRPOINTER_REG_2__SCAN_IN : (~P2_PHYADDRPOINTER_REG_1__SCAN_IN ^ P2_PHYADDRPOINTER_REG_2__SCAN_IN)));
  assign new_n4127_ = new_n4096_ & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_));
  assign new_n4128_ = new_n4129_ & new_n4169_ & new_n4141_ & new_n4150_ & ~new_n4185_ & new_n4176_ & new_n4182_;
  assign new_n4129_ = new_n4130_ & ((~new_n4132_ & P2_INSTQUEUE_REG_0__1__SCAN_IN) | new_n4136_ | ~new_n4139_) & (~new_n4140_ | (~new_n3097_ & P1_INSTQUEUE_REG_9__7__SCAN_IN));
  assign new_n4130_ = (~new_n3007_ | (~new_n3038_ & (~new_n3036_ | (~new_n3035_ & P1_STATEBS16_REG_SCAN_IN)))) & (new_n4131_ | (~new_n3044_ & new_n3047_));
  assign new_n4131_ = ~P1_INSTQUEUE_REG_3__0__SCAN_IN & ~P1_INSTQUEUE_REG_3__3__SCAN_IN;
  assign new_n4132_ = new_n4135_ & ((~new_n2969_ & (~new_n4133_ | ~new_n2968_)) | ((~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ (P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & (~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | (P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & (P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)));
  assign new_n4133_ = (~new_n4134_ | ~new_n1670_ | (new_n1664_ & (~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_))) | (~new_n1664_ & ((new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_)))) | (~new_n1412_ & (new_n1409_ | ~new_n1421_) & (~new_n1409_ | new_n1421_)) | (new_n1412_ & (new_n1409_ ^ new_n1421_))) & (new_n1670_ | new_n1666_ | (new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) | (~new_n1412_ ^ (~new_n1409_ ^ new_n1421_)));
  assign new_n4134_ = (new_n1315_ & P2_INSTQUEUE_REG_0__1__SCAN_IN) ^ (~new_n1417_ | (new_n1413_ & new_n1407_));
  assign new_n4135_ = new_n2966_ & (new_n3537_ | (~P2_STATE2_REG_3__SCAN_IN & (new_n1809_ | ~P2_STATE2_REG_2__SCAN_IN)));
  assign new_n4136_ = new_n3115_ & (new_n4137_ | (new_n4138_ & (new_n4133_ | ~P2_STATEBS16_REG_SCAN_IN)));
  assign new_n4137_ = P2_STATE2_REG_2__SCAN_IN & (new_n1809_ | new_n3537_);
  assign new_n4138_ = new_n2970_ & (~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ (P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & (~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | (P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & (P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  assign new_n4139_ = (~new_n3199_ | ~new_n3244_) & (~new_n3187_ | ~new_n3241_) & (~new_n3537_ | new_n1322_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n4140_ = (~new_n3049_ | new_n3106_) & (~new_n3031_ | ~new_n3124_) & (~new_n3103_ | ~new_n3155_) & (~new_n4068_ | ~new_n3100_);
  assign new_n4141_ = (new_n4143_ | ~new_n4144_ | (~new_n3389_ & P2_INSTQUEUE_REG_3__7__SCAN_IN)) & (~new_n4148_ | (new_n4142_ & new_n2683_ & ~new_n1335_));
  assign new_n4142_ = (new_n1312_ & new_n1315_ & P2_INSTQUEUE_REG_0__7__SCAN_IN) ? new_n1443_ : (new_n1315_ & ~new_n1443_);
  assign new_n4143_ = new_n3113_ & ((P2_STATE2_REG_2__SCAN_IN & (new_n1808_ | new_n3370_)) | ((~new_n3369_ | ~P2_STATEBS16_REG_SCAN_IN) & new_n3371_ & ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN));
  assign new_n4144_ = (~new_n4145_ | ~new_n4083_) & ~new_n4147_ & (~new_n4146_ | ~new_n2968_ | ~new_n3274_);
  assign new_n4145_ = ~new_n1670_ & new_n1666_ & (~new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ ^ (~new_n1409_ ^ new_n1421_));
  assign new_n4146_ = new_n3059_ & (~new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ ^ (~new_n1409_ ^ new_n1421_));
  assign new_n4147_ = new_n3370_ & ~new_n1335_ & new_n2966_ & P2_STATE2_REG_3__SCAN_IN;
  assign new_n4148_ = (~new_n4149_ | ~new_n2683_ | ~new_n1335_) & (new_n2683_ | ~P2_EBX_REG_8__SCAN_IN);
  assign new_n4149_ = ~new_n1985_ ^ (new_n1978_ & ~new_n1984_);
  assign new_n4150_ = (new_n4151_ ? (P2_STATE2_REG_2__SCAN_IN & P2_STATE2_REG_1__SCAN_IN) : (P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN)) & (new_n4167_ | ~new_n4168_ | (~new_n3246_ & P2_INSTQUEUE_REG_13__6__SCAN_IN));
  assign new_n4151_ = P2_STATE2_REG_0__SCAN_IN & (~new_n4166_ | (P2_STATE2_REG_0__SCAN_IN & (~new_n4163_ | (~new_n4152_ & new_n4160_))));
  assign new_n4152_ = (P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | (~new_n4153_ & ~new_n4154_)) & (new_n4156_ | P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) & ((new_n4156_ & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN) | (new_n4157_ & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (new_n4159_ & (new_n4157_ | P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)));
  assign new_n4153_ = P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~new_n3177_ & new_n3178_;
  assign new_n4154_ = (new_n3177_ | ~new_n3178_) & (~new_n4155_ | (~new_n3171_ & (~new_n1327_ | (~new_n1383_ & (new_n1386_ | new_n1387_))) & (new_n1327_ | new_n1383_ | (~new_n1386_ & ~new_n1387_))));
  assign new_n4155_ = (new_n3174_ | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) | (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN))) & (new_n3255_ | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) | (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN & (~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN))) & (~new_n3254_ | (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) | ((~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN) & (P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN)));
  assign new_n4156_ = (~new_n3177_ & new_n3178_) ? ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN : (new_n3253_ & (new_n3171_ | (new_n1387_ & ~new_n1410_) | (~new_n1387_ & new_n1410_)));
  assign new_n4157_ = (~new_n3177_ & new_n3178_) ? ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN : (new_n4158_ & (~new_n1413_ | new_n3171_));
  assign new_n4158_ = (new_n3174_ | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (new_n3175_ | ~new_n1367_ | (P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN));
  assign new_n4159_ = (~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | new_n3177_ | ~new_n3178_) & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & (new_n3170_ | (~new_n3177_ & new_n3178_));
  assign new_n4160_ = (new_n4161_ | ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN) & (~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | new_n4153_ | new_n4154_);
  assign new_n4161_ = (~new_n3177_ & new_n3178_) ? P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN : (new_n1786_ & new_n1322_ & (~new_n4162_ | new_n1367_ | ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN) & (new_n4162_ | (~new_n1367_ & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN)));
  assign new_n4162_ = P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign new_n4163_ = ~new_n4161_ & new_n4164_ & (new_n4156_ | (~new_n4153_ & ~new_n4154_));
  assign new_n4164_ = (~new_n3554_ | (~P2_FLUSH_REG_SCAN_IN & ~P2_MORE_REG_SCAN_IN)) & (new_n3169_ | (~new_n1783_ & ~new_n2667_)) & new_n4165_ & (~new_n3169_ | ~new_n2684_);
  assign new_n4165_ = (new_n2668_ | new_n1788_) & ~P2_STATE2_REG_1__SCAN_IN & (~new_n2708_ | new_n1370_);
  assign new_n4166_ = (~new_n1376_ | P2_STATE_REG_0__SCAN_IN | new_n1790_ | P2_STATEBS16_REG_SCAN_IN) & P2_STATE2_REG_2__SCAN_IN & (P2_STATE2_REG_0__SCAN_IN | (new_n1790_ & P2_STATE2_REG_1__SCAN_IN));
  assign new_n4167_ = new_n3191_ & ((P2_STATE2_REG_2__SCAN_IN & (new_n1806_ | (new_n3063_ & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN))) | ((~new_n3159_ | ~P2_STATEBS16_REG_SCAN_IN) & new_n3063_ & ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN));
  assign new_n4168_ = (~new_n3060_ | ~new_n3193_) & (~new_n3081_ | ~new_n3195_) & (~new_n3248_ | new_n1317_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n4169_ = new_n4170_ & (new_n4172_ | ~new_n4173_ | (~new_n3389_ & P2_INSTQUEUE_REG_3__1__SCAN_IN)) & (new_n4174_ | ~new_n4175_ | (~new_n3389_ & P2_INSTQUEUE_REG_3__6__SCAN_IN));
  assign new_n4170_ = ~new_n4171_ & (~new_n2982_ | (~new_n3066_ & (~new_n3067_ | (P2_STATEBS16_REG_SCAN_IN & (new_n3058_ | new_n3060_)))));
  assign new_n4171_ = new_n3155_ & (new_n2994_ ? ((new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ | (~new_n2148_ & ~new_n2200_) | (new_n2148_ & new_n2200_)) & (~new_n2154_ | (~new_n2148_ ^ ~new_n2200_))) : (new_n2284_ & (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & (new_n2154_ ^ (~new_n2148_ ^ ~new_n2200_))));
  assign new_n4172_ = new_n3115_ & ((P2_STATE2_REG_2__SCAN_IN & (new_n1808_ | new_n3370_)) | ((~new_n3369_ | ~P2_STATEBS16_REG_SCAN_IN) & new_n3371_ & ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN));
  assign new_n4173_ = (~new_n4145_ | ~new_n3241_) & (~new_n4146_ | ~new_n3244_) & (~new_n3370_ | new_n1322_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n4174_ = new_n3191_ & ((P2_STATE2_REG_2__SCAN_IN & (new_n1808_ | new_n3370_)) | ((~new_n3369_ | ~P2_STATEBS16_REG_SCAN_IN) & new_n3371_ & ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN));
  assign new_n4175_ = (~new_n4145_ | ~new_n3193_) & (~new_n4146_ | ~new_n3195_) & (~new_n3370_ | new_n1317_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n4176_ = (new_n4179_ | ~P2_INSTQUEUE_REG_10__6__SCAN_IN) & ((~new_n3246_ & P2_INSTQUEUE_REG_13__7__SCAN_IN) | ~new_n4177_ | (~new_n3158_ & new_n3113_));
  assign new_n4177_ = (~new_n3060_ | ~new_n4083_) & ~new_n4178_ & (~new_n3081_ | ~new_n2968_ | ~new_n3274_);
  assign new_n4178_ = new_n3248_ & ~new_n1335_ & new_n2966_ & P2_STATE2_REG_3__SCAN_IN;
  assign new_n4179_ = new_n4181_ & ((~new_n1418_ & new_n3364_) | (~new_n2969_ & (new_n4180_ | ~new_n2968_)));
  assign new_n4180_ = ~new_n3242_ & ~new_n3059_ & (~new_n1664_ | (new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_))) & (new_n1664_ | ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ ^ (~new_n1409_ ^ new_n1421_));
  assign new_n4181_ = new_n2966_ & (new_n3538_ | (~P2_STATE2_REG_3__SCAN_IN & (new_n1802_ | ~P2_STATE2_REG_2__SCAN_IN)));
  assign new_n4182_ = (~new_n1686_ | (~new_n2665_ & ~new_n2678_)) & ((~new_n3246_ & P2_INSTQUEUE_REG_13__0__SCAN_IN) | ~new_n4183_ | (~new_n3158_ & new_n2982_));
  assign new_n4183_ = (~new_n3060_ | ~new_n2968_ | ~new_n2981_) & ~new_n4184_ & (~new_n3081_ | ~new_n2968_ | ~new_n2975_);
  assign new_n4184_ = new_n3248_ & ~new_n1370_ & new_n2966_ & P2_STATE2_REG_3__SCAN_IN;
  assign new_n4185_ = new_n2004_ & (new_n3402_ | (~new_n1995_ ^ (~new_n1994_ & new_n1977_ & ~new_n1993_)));
  assign new_n4186_ = new_n4187_ & new_n4198_ & new_n4209_ & new_n4221_ & new_n4223_ & ~new_n4236_ & (new_n4233_ | ~P1_INSTQUEUE_REG_10__7__SCAN_IN);
  assign new_n4187_ = (new_n4188_ | ~new_n4191_ | (~new_n3039_ & new_n4197_)) & (new_n4192_ | ~new_n4195_ | (~new_n3029_ & new_n3049_));
  assign new_n4188_ = P1_INSTQUEUE_REG_6__0__SCAN_IN & (~new_n4190_ | (new_n3041_ & ~new_n4189_));
  assign new_n4189_ = ~new_n2998_ & (~new_n2996_ | (new_n2994_ & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ | (~new_n2148_ & ~new_n2200_) | (new_n2148_ & new_n2200_)) & (~new_n2154_ | (~new_n2148_ ^ ~new_n2200_))) | (~new_n2994_ & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & new_n2284_ & (new_n2154_ | (~new_n2148_ & ~new_n2200_) | (new_n2148_ & new_n2200_)) & (~new_n2154_ | (~new_n2148_ ^ ~new_n2200_))));
  assign new_n4190_ = new_n3003_ & (~P1_STATE2_REG_3__SCAN_IN | (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN)) & (~P1_STATE2_REG_2__SCAN_IN | (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)));
  assign new_n4191_ = (~new_n3265_ | ~new_n2996_ | new_n3230_) & (~new_n3352_ | ~new_n3042_) & (~new_n3266_ | ~new_n2996_ | new_n3123_);
  assign new_n4192_ = P1_INSTQUEUE_REG_8__7__SCAN_IN & (~new_n4194_ | (new_n3032_ & ~new_n4193_));
  assign new_n4193_ = ~new_n2998_ & (~new_n2996_ | (~new_n2994_ & (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ ^ (~new_n2148_ ^ ~new_n2200_))) | (new_n2994_ & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & new_n2284_ & (new_n2154_ | (~new_n2148_ & ~new_n2200_) | (new_n2148_ & new_n2200_)) & (~new_n2154_ | (~new_n2148_ ^ ~new_n2200_))));
  assign new_n4194_ = new_n3003_ & (~P1_STATE2_REG_2__SCAN_IN | ((P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ^ (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)) & (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ^ ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)))) & (~P1_STATE2_REG_3__SCAN_IN | (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN));
  assign new_n4195_ = (~new_n3030_ | ~new_n3124_) & ~new_n4196_ & (~new_n3031_ | ~new_n3155_);
  assign new_n4196_ = new_n4068_ & ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n4197_ = new_n3003_ & (new_n2954_ ? BUF1_REG_0__SCAN_IN : DATAI_0_);
  assign new_n4198_ = ~new_n4201_ & (~new_n4199_ | (~new_n3034_ & new_n3053_) | (P1_INSTQUEUE_REG_4__5__SCAN_IN & (~new_n4208_ | (new_n4206_ & ~new_n4207_))));
  assign new_n4199_ = ~new_n4200_ & (~new_n3152_ | ~new_n3055_) & (~new_n3056_ | ~new_n3037_);
  assign new_n4200_ = new_n3054_ & new_n2284_ & new_n2994_ & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & (new_n2154_ ^ (~new_n2148_ ^ ~new_n2200_));
  assign new_n4201_ = (~new_n2937_ | (~new_n4202_ & new_n4203_)) & (~P3_INSTADDRPOINTER_REG_22__SCAN_IN | new_n2937_ | new_n3282_) & (~P3_REIP_REG_22__SCAN_IN | P3_STATE2_REG_2__SCAN_IN | (~new_n2937_ & ~new_n3282_));
  assign new_n4202_ = ((new_n2925_ ^ ~P3_INSTADDRPOINTER_REG_22__SCAN_IN) | new_n2930_ | (~new_n2925_ & ~new_n2936_)) & new_n2935_ & ((new_n2925_ & ~P3_INSTADDRPOINTER_REG_22__SCAN_IN) | (~new_n2925_ & P3_INSTADDRPOINTER_REG_22__SCAN_IN) | (~new_n2930_ & (new_n2925_ | new_n2936_)));
  assign new_n4203_ = ((~new_n2864_ & ~P3_INSTADDRPOINTER_REG_22__SCAN_IN) | ~new_n2928_ | (new_n2864_ & P3_INSTADDRPOINTER_REG_22__SCAN_IN)) & new_n4204_ & ((~new_n2912_ & ~P3_INSTADDRPOINTER_REG_22__SCAN_IN) | ~new_n2926_ | (new_n2912_ & P3_INSTADDRPOINTER_REG_22__SCAN_IN));
  assign new_n4204_ = (new_n4205_ | (P3_INSTADDRPOINTER_REG_22__SCAN_IN & new_n2843_ & new_n2786_) | (~P3_INSTADDRPOINTER_REG_22__SCAN_IN & (~new_n2843_ | ~new_n2786_))) & (new_n3287_ | (P3_INSTADDRPOINTER_REG_22__SCAN_IN & new_n2780_ & new_n2786_) | (~P3_INSTADDRPOINTER_REG_22__SCAN_IN & (~new_n2780_ | ~new_n2786_))) & (~new_n2850_ | (P3_INSTADDRPOINTER_REG_22__SCAN_IN & new_n2848_ & new_n2786_) | (~P3_INSTADDRPOINTER_REG_22__SCAN_IN & (~new_n2848_ | ~new_n2786_)));
  assign new_n4205_ = (~new_n2846_ | ~new_n2809_) & new_n2857_ & ~new_n2858_ & ~new_n2859_ & new_n2860_ & (~new_n2846_ | new_n2809_);
  assign new_n4206_ = ~new_n3037_ & (~new_n2990_ | ~new_n2133_ | ~new_n2986_ | new_n2987_);
  assign new_n4207_ = ~new_n2998_ & (~new_n2996_ | (new_n2284_ & new_n2994_ & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & (new_n2154_ ^ (~new_n2148_ ^ ~new_n2200_))) | (~new_n2994_ & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & ~new_n2284_ & (new_n2154_ | (~new_n2148_ & ~new_n2200_) | (new_n2148_ & new_n2200_)) & (~new_n2154_ | (~new_n2148_ ^ ~new_n2200_))));
  assign new_n4208_ = new_n3003_ & (~P1_STATE2_REG_2__SCAN_IN | (~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ^ ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)))) & (~P1_STATE2_REG_3__SCAN_IN | (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN));
  assign new_n4209_ = (new_n4211_ | new_n4212_) & (new_n4217_ | (~new_n3007_ & ~new_n3049_)) & (~new_n4215_ | (~new_n4210_ & P1_INSTQUEUE_REG_15__2__SCAN_IN));
  assign new_n4210_ = new_n3259_ & (~new_n3258_ | (~new_n2998_ & (~new_n2996_ | (new_n2276_ & new_n3257_))));
  assign new_n4211_ = ~new_n3053_ & ~new_n4197_;
  assign new_n4212_ = ~new_n4214_ & ((~new_n4213_ & P1_STATEBS16_REG_SCAN_IN) | ~new_n2576_ | (~new_n3353_ & (~new_n2985_ | ~new_n2990_ | new_n2133_)));
  assign new_n4213_ = new_n2994_ ? ((~new_n2277_ & (new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_))) | (new_n2277_ & ((~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_)))) | new_n2284_ | (~new_n2154_ & (~new_n2148_ | ~new_n2200_) & (new_n2148_ | new_n2200_)) | (new_n2154_ & (~new_n2148_ ^ new_n2200_))) : ((~new_n2277_ & (new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_))) | (new_n2277_ & ((~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_)))) | ~new_n2284_ | (~new_n2154_ & (~new_n2148_ | ~new_n2200_) & (new_n2148_ | new_n2200_)) | (new_n2154_ & (~new_n2148_ ^ new_n2200_)));
  assign new_n4214_ = P1_STATE2_REG_2__SCAN_IN & new_n2120_ & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n4215_ = (~new_n3024_ | new_n3221_) & (~new_n3121_ | ~new_n3026_) & ~new_n4216_ & (~new_n4098_ | ~new_n3027_);
  assign new_n4216_ = new_n3223_ & ~new_n2097_ & new_n3003_ & P1_STATE2_REG_3__SCAN_IN;
  assign new_n4217_ = ~new_n4220_ & (new_n4218_ | ~new_n2576_ | (P1_STATEBS16_REG_SCAN_IN & (new_n3161_ | new_n4098_)));
  assign new_n4218_ = ~new_n4219_ & (new_n2989_ | new_n2990_ | ~new_n2986_ | new_n2987_);
  assign new_n4219_ = ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n4220_ = P1_STATE2_REG_2__SCAN_IN & (P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)) & (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ^ P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN));
  assign new_n4221_ = (~new_n4222_ | (~new_n4210_ & P1_INSTQUEUE_REG_15__7__SCAN_IN)) & (~new_n2665_ | (~new_n1644_ & new_n1620_) | (new_n1644_ & ~new_n1620_));
  assign new_n4222_ = (~new_n3049_ | new_n3221_) & (~new_n3121_ | ~new_n3124_) & (~new_n4098_ | ~new_n3155_) & (~new_n4068_ | ~new_n3223_);
  assign new_n4223_ = (~new_n4227_ | (~new_n4224_ & P1_INSTQUEUE_REG_13__3__SCAN_IN)) & (new_n4231_ | ~new_n4232_ | (~new_n4229_ & P1_INSTQUEUE_REG_1__7__SCAN_IN));
  assign new_n4224_ = new_n4226_ & (~new_n4225_ | (~new_n2998_ & (new_n3378_ | ~new_n2996_)));
  assign new_n4225_ = ~new_n3214_ & (~new_n3004_ | ~new_n2990_ | new_n2133_);
  assign new_n4226_ = new_n3003_ & ((~P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_2__SCAN_IN) | ((P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_STATE2_REG_3__SCAN_IN) & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN));
  assign new_n4227_ = (~new_n3109_ | new_n3212_) & (~new_n3104_ | ~new_n3378_ | new_n2994_) & ~new_n4228_ & (~new_n3105_ | ~new_n3378_ | ~new_n2994_);
  assign new_n4228_ = new_n3214_ & ~new_n2091_ & new_n3003_ & P1_STATE2_REG_3__SCAN_IN;
  assign new_n4229_ = new_n4230_ & (new_n3219_ | (new_n2988_ & new_n3004_) | (~new_n2998_ & (new_n3217_ | ~new_n2996_)));
  assign new_n4230_ = new_n3003_ & (new_n3219_ | (~P1_STATE2_REG_3__SCAN_IN & (new_n4219_ | ~P1_STATE2_REG_2__SCAN_IN)));
  assign new_n4231_ = new_n3049_ & (new_n3218_ | ((~new_n3217_ | ~P1_STATEBS16_REG_SCAN_IN) & new_n2576_ & (new_n3219_ | (new_n2988_ & new_n3004_))));
  assign new_n4232_ = (~new_n3161_ | ~new_n3124_) & (~new_n4068_ | ~new_n3219_) & (~new_n2993_ | ~new_n3155_);
  assign new_n4233_ = new_n4234_ & (new_n4235_ | (new_n2985_ & new_n3092_) | (~new_n2998_ & (~new_n2996_ | new_n3103_ | new_n3397_)));
  assign new_n4234_ = new_n3003_ & (~P1_STATE2_REG_3__SCAN_IN | (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN)) & (~P1_STATE2_REG_2__SCAN_IN | (~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)));
  assign new_n4235_ = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n4236_ = ((new_n2269_ & new_n2271_) | (~new_n2269_ & ~new_n2271_) | ((~new_n2282_ | (new_n2278_ & (~new_n2276_ | ~new_n2237_))) & (new_n2278_ | ~new_n2276_ | ~new_n2237_))) & ~new_n2630_ & ~new_n3386_ & ((new_n2269_ ^ new_n2271_) | (new_n2282_ & (~new_n2278_ | (new_n2276_ & new_n2237_))) | (~new_n2278_ & new_n2276_ & new_n2237_));
  assign new_n4237_ = new_n4238_ & new_n4327_ & new_n4264_ & new_n4284_ & new_n4292_ & new_n4317_ & new_n4299_ & new_n4308_;
  assign new_n4238_ = ~new_n4239_ & ~new_n4245_ & (~new_n4249_ | (~new_n3091_ & P1_INSTQUEUE_REG_11__7__SCAN_IN)) & ~new_n4255_ & (~new_n4261_ | (~new_n3091_ & P1_INSTQUEUE_REG_11__2__SCAN_IN));
  assign new_n4239_ = (new_n4240_ | ~new_n2937_) & (~P3_INSTADDRPOINTER_REG_19__SCAN_IN | new_n2937_ | new_n3282_) & (~P3_REIP_REG_19__SCAN_IN | P3_STATE2_REG_2__SCAN_IN | (~new_n2937_ & ~new_n3282_));
  assign new_n4240_ = new_n4242_ & (((new_n4241_ | ~P3_INSTADDRPOINTER_REG_19__SCAN_IN) & (~new_n2923_ | new_n2906_) & (~new_n4241_ | P3_INSTADDRPOINTER_REG_19__SCAN_IN)) | ~new_n2927_ | new_n2906_ | (new_n2923_ & (new_n4241_ ^ P3_INSTADDRPOINTER_REG_19__SCAN_IN)));
  assign new_n4241_ = (new_n2925_ | ~P3_INSTADDRPOINTER_REG_18__SCAN_IN) & (new_n2925_ | (~P3_INSTADDRPOINTER_REG_17__SCAN_IN & ~P3_INSTADDRPOINTER_REG_16__SCAN_IN & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_15__SCAN_IN) & ((new_n2925_ & ~P3_INSTADDRPOINTER_REG_15__SCAN_IN) | ((new_n2925_ | ~P3_INSTADDRPOINTER_REG_14__SCAN_IN) & (new_n2931_ | (new_n2925_ & ~P3_INSTADDRPOINTER_REG_14__SCAN_IN)))))) & ((new_n2925_ & ~P3_INSTADDRPOINTER_REG_15__SCAN_IN) | ((new_n2925_ | ~P3_INSTADDRPOINTER_REG_14__SCAN_IN) & (new_n2931_ | (new_n2925_ & ~P3_INSTADDRPOINTER_REG_14__SCAN_IN))) | ~P3_INSTADDRPOINTER_REG_17__SCAN_IN | ~P3_INSTADDRPOINTER_REG_16__SCAN_IN | ~P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  assign new_n4242_ = ~new_n4243_ & new_n4244_ & (~new_n2928_ | (new_n3357_ & P3_INSTADDRPOINTER_REG_19__SCAN_IN) | (~new_n3357_ & ~P3_INSTADDRPOINTER_REG_19__SCAN_IN));
  assign new_n4243_ = (P3_INSTADDRPOINTER_REG_19__SCAN_IN | (new_n2781_ & new_n2924_ & (new_n2913_ | ~new_n2922_))) & new_n2926_ & (~P3_INSTADDRPOINTER_REG_19__SCAN_IN | ~new_n2781_ | ~new_n2924_ | (~new_n2913_ & new_n2922_));
  assign new_n4244_ = (new_n4205_ | (~new_n2843_ & ~P3_INSTADDRPOINTER_REG_19__SCAN_IN) | (P3_INSTADDRPOINTER_REG_0__SCAN_IN & new_n2780_ & P3_INSTADDRPOINTER_REG_19__SCAN_IN)) & (~new_n2850_ | (new_n2848_ & P3_INSTADDRPOINTER_REG_19__SCAN_IN) | (~new_n2848_ & ~P3_INSTADDRPOINTER_REG_19__SCAN_IN)) & (new_n3287_ | (~new_n2780_ & ~P3_INSTADDRPOINTER_REG_19__SCAN_IN) | (new_n2780_ & P3_INSTADDRPOINTER_REG_19__SCAN_IN));
  assign new_n4245_ = (new_n4246_ | ~new_n2937_) & (~P3_INSTADDRPOINTER_REG_20__SCAN_IN | new_n2937_ | new_n3282_) & (~P3_REIP_REG_20__SCAN_IN | P3_STATE2_REG_2__SCAN_IN | (~new_n2937_ & ~new_n3282_));
  assign new_n4246_ = (~new_n2935_ | (((new_n2925_ & (new_n4241_ | ~P3_INSTADDRPOINTER_REG_19__SCAN_IN)) | (new_n4241_ & ~P3_INSTADDRPOINTER_REG_19__SCAN_IN) | (new_n2925_ & P3_INSTADDRPOINTER_REG_20__SCAN_IN) | (~new_n2925_ & ~P3_INSTADDRPOINTER_REG_20__SCAN_IN)) & ((~new_n2925_ & (~new_n4241_ | P3_INSTADDRPOINTER_REG_19__SCAN_IN)) | (~new_n4241_ & P3_INSTADDRPOINTER_REG_19__SCAN_IN) | (new_n2925_ ^ P3_INSTADDRPOINTER_REG_20__SCAN_IN)))) & new_n4247_ & ((~P3_INSTADDRPOINTER_REG_20__SCAN_IN & (~new_n3357_ | ~P3_INSTADDRPOINTER_REG_19__SCAN_IN)) | ~new_n2928_ | (new_n3357_ & P3_INSTADDRPOINTER_REG_19__SCAN_IN & P3_INSTADDRPOINTER_REG_20__SCAN_IN));
  assign new_n4247_ = new_n4248_ & ((~P3_INSTADDRPOINTER_REG_20__SCAN_IN & (~P3_INSTADDRPOINTER_REG_19__SCAN_IN | ~new_n2781_ | ~new_n2924_ | (~new_n2913_ & new_n2922_))) | ~new_n2926_ | (P3_INSTADDRPOINTER_REG_20__SCAN_IN & P3_INSTADDRPOINTER_REG_19__SCAN_IN & new_n2781_ & new_n2924_ & (new_n2913_ | ~new_n2922_)));
  assign new_n4248_ = (new_n4205_ | (~P3_INSTADDRPOINTER_REG_20__SCAN_IN & (~P3_INSTADDRPOINTER_REG_0__SCAN_IN | ~new_n2780_ | ~P3_INSTADDRPOINTER_REG_19__SCAN_IN)) | (P3_INSTADDRPOINTER_REG_20__SCAN_IN & P3_INSTADDRPOINTER_REG_0__SCAN_IN & new_n2780_ & P3_INSTADDRPOINTER_REG_19__SCAN_IN)) & (~new_n2850_ | (P3_INSTADDRPOINTER_REG_20__SCAN_IN & new_n2848_ & P3_INSTADDRPOINTER_REG_19__SCAN_IN) | (~P3_INSTADDRPOINTER_REG_20__SCAN_IN & (~new_n2848_ | ~P3_INSTADDRPOINTER_REG_19__SCAN_IN))) & (new_n3287_ | (P3_INSTADDRPOINTER_REG_20__SCAN_IN & new_n2780_ & P3_INSTADDRPOINTER_REG_19__SCAN_IN) | (~P3_INSTADDRPOINTER_REG_20__SCAN_IN & (~new_n2780_ | ~P3_INSTADDRPOINTER_REG_19__SCAN_IN)));
  assign new_n4249_ = (~new_n3049_ | new_n4250_) & new_n4253_ & (~new_n3397_ | ~new_n3124_);
  assign new_n4250_ = ~new_n4252_ & (~new_n4251_ | (P1_STATEBS16_REG_SCAN_IN & new_n2284_ & (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & (new_n2154_ ^ (new_n2148_ ^ new_n2200_))));
  assign new_n4251_ = new_n2576_ & (new_n3095_ | (new_n2987_ & (~new_n2050_ | ~new_n2143_) & (new_n2050_ | new_n2143_) & (new_n2133_ | new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_)))) & (~new_n2133_ | (~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_))))) & (new_n2131_ ^ ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_))))));
  assign new_n4252_ = P1_STATE2_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n4253_ = ~new_n4254_ & (~new_n3155_ | ~new_n2284_ | ~new_n2994_ | (~new_n2277_ & (new_n2154_ | (new_n2148_ & new_n2200_)) & (new_n2148_ | new_n2200_)) | (new_n2277_ & ((~new_n2154_ & (~new_n2148_ | ~new_n2200_)) | (~new_n2148_ & ~new_n2200_))) | (~new_n2154_ ^ (new_n2148_ ^ new_n2200_)));
  assign new_n4254_ = new_n4068_ & new_n3095_;
  assign new_n4255_ = (~P1_INSTQUEUE_REG_3__5__SCAN_IN | (~new_n3044_ & new_n3047_)) & (~new_n3053_ | new_n4256_) & new_n4259_ & (~new_n2995_ | ~new_n3054_);
  assign new_n4256_ = ~new_n4258_ & (~new_n4257_ | (P1_STATEBS16_REG_SCAN_IN & new_n2284_ & (new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & (new_n2154_ ^ (new_n2148_ ^ new_n2200_))));
  assign new_n4257_ = new_n2576_ & (new_n3046_ | (new_n2987_ & (~new_n2050_ | ~new_n2143_) & (new_n2050_ | new_n2143_) & (new_n2133_ ^ (~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_))))) & (new_n2131_ ^ ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_))))));
  assign new_n4258_ = P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & new_n2992_ & P1_STATE2_REG_2__SCAN_IN;
  assign new_n4259_ = ~new_n4260_ & (~new_n3055_ | ~new_n2284_ | ~new_n2994_ | (~new_n2277_ ^ ((new_n2154_ | (new_n2148_ & new_n2200_)) & (new_n2148_ | new_n2200_))) | (~new_n2154_ ^ (new_n2148_ ^ new_n2200_)));
  assign new_n4260_ = new_n3056_ & new_n3046_;
  assign new_n4261_ = (~new_n3024_ | new_n4250_) & new_n4262_ & (~new_n3397_ | ~new_n3026_);
  assign new_n4262_ = ~new_n4263_ & (~new_n3027_ | ~new_n2284_ | ~new_n2994_ | (~new_n2277_ & (new_n2154_ | (new_n2148_ & new_n2200_)) & (new_n2148_ | new_n2200_)) | (new_n2277_ & ((~new_n2154_ & (~new_n2148_ | ~new_n2200_)) | (~new_n2148_ & ~new_n2200_))) | (~new_n2154_ ^ (new_n2148_ ^ new_n2200_)));
  assign new_n4263_ = new_n3095_ & ~new_n2097_ & P1_STATE2_REG_3__SCAN_IN & ~P1_STATE2_REG_0__SCAN_IN & (new_n2997_ | (~new_n2477_ & P1_STATE2_REG_3__SCAN_IN));
  assign new_n4264_ = (~new_n4268_ | (~new_n4265_ & P2_INSTQUEUE_REG_9__6__SCAN_IN)) & ~new_n4279_ & ~new_n4283_ & ~new_n4275_ & (new_n4229_ | ~P1_INSTQUEUE_REG_1__5__SCAN_IN);
  assign new_n4265_ = new_n4267_ & ((new_n3364_ & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) | (~new_n2969_ & (~new_n4266_ | ~new_n2968_)));
  assign new_n4266_ = (new_n4134_ | ~new_n1670_ | (new_n1664_ & (~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_))) | (~new_n1664_ & ((new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_)))) | (~new_n1412_ ^ (~new_n1409_ ^ new_n1421_))) & (new_n1666_ | new_n1670_ | ((new_n4134_ & new_n1670_) ? ((new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) | (~new_n1412_ & (new_n1409_ | ~new_n1421_) & (~new_n1409_ | new_n1421_)) | (new_n1412_ & (new_n1409_ ^ new_n1421_))) : ((new_n1664_ & (~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_))) | (~new_n1664_ & ((new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_)))) | (~new_n1412_ ^ (~new_n1409_ ^ new_n1421_)))));
  assign new_n4267_ = new_n2966_ & ((~P2_STATE2_REG_3__SCAN_IN & (new_n1819_ | ~P2_STATE2_REG_2__SCAN_IN)) | (new_n3364_ & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN));
  assign new_n4268_ = new_n4272_ & (~new_n4270_ | ~new_n3193_) & (~new_n3191_ | (~new_n4271_ & (~new_n4274_ | (P2_STATEBS16_REG_SCAN_IN & (new_n4269_ | new_n4270_)))));
  assign new_n4269_ = new_n2963_ & (~new_n1664_ | (new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_))) & (new_n1664_ | ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ ^ (~new_n1409_ ^ new_n1421_));
  assign new_n4270_ = new_n3242_ & (new_n3059_ ? ((~new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ | (~new_n1409_ & new_n1421_) | (new_n1409_ & ~new_n1421_)) & (~new_n1412_ | (~new_n1409_ ^ new_n1421_))) : ((~new_n1664_ | (new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_))) & (new_n1664_ | ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) & (new_n1412_ ^ (~new_n1409_ ^ new_n1421_))));
  assign new_n4271_ = P2_STATE2_REG_2__SCAN_IN & (new_n1819_ | (new_n3364_ & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN));
  assign new_n4272_ = ~new_n4273_ & (~new_n3195_ | ~new_n2963_ | (new_n1664_ & (~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_))) | (~new_n1664_ & ((new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_)))) | (~new_n1412_ ^ (new_n1409_ ^ ~new_n1421_)));
  assign new_n4273_ = ~new_n1317_ & new_n2966_ & P2_STATE2_REG_3__SCAN_IN & new_n3364_ & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n4274_ = new_n2970_ & new_n3364_ & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n4275_ = ~new_n4278_ & ((~P2_STATE2_REG_0__SCAN_IN & (new_n4276_ | (new_n4166_ & (~P2_STATE2_REG_0__SCAN_IN | (new_n4163_ & (new_n4152_ | ~new_n4160_)))))) | (P2_STATE2_REG_0__SCAN_IN & (~new_n4166_ | (P2_STATE2_REG_0__SCAN_IN & (~new_n4163_ | (~new_n4152_ & new_n4160_)))) & (~new_n4277_ | (new_n4163_ & (new_n4152_ | ~new_n4160_)))));
  assign new_n4276_ = new_n2022_ & new_n3169_ & P2_STATE2_REG_3__SCAN_IN;
  assign new_n4277_ = P2_STATE2_REG_2__SCAN_IN & (new_n2011_ | ~P2_STATE2_REG_1__SCAN_IN);
  assign new_n4278_ = ~P2_STATE2_REG_2__SCAN_IN & P2_STATE2_REG_0__SCAN_IN & (new_n1790_ | (P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_1__SCAN_IN));
  assign new_n4279_ = new_n3191_ & (new_n4280_ | new_n4281_ | new_n4137_ | (new_n4138_ & (new_n4133_ | ~P2_STATEBS16_REG_SCAN_IN)));
  assign new_n4280_ = P2_STATE2_REG_2__SCAN_IN & (new_n1802_ | new_n3538_);
  assign new_n4281_ = new_n4282_ & (~P2_STATEBS16_REG_SCAN_IN | new_n3242_ | new_n3059_ | (new_n1664_ & (~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_))) | (~new_n1664_ & ((new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_)))) | (~new_n1412_ ^ (~new_n1409_ ^ new_n1421_)));
  assign new_n4282_ = new_n2970_ & ~new_n1418_ & new_n3364_;
  assign new_n4283_ = P2_INSTQUEUE_REG_12__0__SCAN_IN & (~new_n3061_ | (~new_n3064_ & (new_n2969_ | (new_n2968_ & ~new_n3058_ & ~new_n3060_))));
  assign new_n4284_ = ((~new_n4265_ & P2_INSTQUEUE_REG_9__1__SCAN_IN) | ~new_n4286_ | (~new_n4285_ & new_n3115_)) & ((~new_n4265_ & P2_INSTQUEUE_REG_9__3__SCAN_IN) | ~new_n4289_ | (~new_n4285_ & new_n3166_));
  assign new_n4285_ = ~new_n4271_ & (~new_n4274_ | (~new_n4266_ & P2_STATEBS16_REG_SCAN_IN));
  assign new_n4286_ = new_n4287_ & (~new_n4270_ | ~new_n3241_);
  assign new_n4287_ = ~new_n4288_ & (~new_n3244_ | ~new_n2963_ | (new_n1664_ & (~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_))) | (~new_n1664_ & ((new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_)))) | (~new_n1412_ ^ (new_n1409_ ^ ~new_n1421_)));
  assign new_n4288_ = ~new_n1322_ & new_n2966_ & P2_STATE2_REG_3__SCAN_IN & new_n3364_ & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n4289_ = new_n4290_ & (~new_n4270_ | ~new_n3211_);
  assign new_n4290_ = ~new_n4291_ & (~new_n2968_ | ~new_n3210_ | ~new_n2963_ | (new_n1664_ & (~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_))) | (~new_n1664_ & ((new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_)))) | (~new_n1412_ ^ (~new_n1409_ ^ new_n1421_)));
  assign new_n4291_ = ~new_n1345_ & new_n2966_ & P2_STATE2_REG_3__SCAN_IN & new_n3364_ & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n4292_ = ~new_n4295_ & ~new_n4296_ & ~new_n4297_ & ~new_n4298_ & new_n4293_ & ~new_n4294_ & (new_n4132_ | ~P2_INSTQUEUE_REG_0__6__SCAN_IN);
  assign new_n4293_ = (new_n4256_ | (~new_n3109_ & ~new_n3049_ & ~new_n4197_)) & (~P1_INSTQUEUE_REG_9__4__SCAN_IN | (~new_n3098_ & new_n3101_));
  assign new_n4294_ = P1_INSTQUEUE_REG_9__1__SCAN_IN & (new_n3098_ | ~new_n3101_);
  assign new_n4295_ = P1_INSTQUEUE_REG_7__4__SCAN_IN & (~new_n3019_ | (new_n3015_ & (new_n2998_ | (~new_n3018_ & new_n2996_))));
  assign new_n4296_ = P2_INSTQUEUE_REG_6__7__SCAN_IN & (~new_n2965_ | ((new_n1418_ | ~new_n2967_) & (new_n2969_ | (new_n2968_ & ~new_n2962_ & ~new_n2964_))));
  assign new_n4297_ = (P2_INSTQUEUE_REG_14__2__SCAN_IN | P2_INSTQUEUE_REG_14__1__SCAN_IN) & (~new_n3083_ | (~new_n3086_ & (new_n2969_ | (new_n2968_ & ~new_n3081_ & ~new_n3082_))));
  assign new_n4298_ = new_n3048_ & ~new_n4250_;
  assign new_n4299_ = ~new_n4307_ & ((~new_n4300_ & P2_INSTQUEUE_REG_4__6__SCAN_IN) | new_n4305_ | ~new_n4306_ | (new_n3393_ & new_n3195_));
  assign new_n4300_ = new_n4302_ & (new_n4304_ | (~new_n2969_ & (~new_n4301_ | ~new_n2968_)));
  assign new_n4301_ = (~new_n3059_ | (new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) | (~new_n1412_ ^ (~new_n1409_ ^ new_n1421_))) & (~new_n3242_ | (new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) | (~new_n1412_ & (new_n1409_ | ~new_n1421_) & (~new_n1409_ | new_n1421_)) | (new_n1412_ & (new_n1409_ ^ new_n1421_)));
  assign new_n4302_ = new_n2966_ & (new_n4303_ | (~P2_STATE2_REG_3__SCAN_IN & (new_n1843_ | ~P2_STATE2_REG_2__SCAN_IN)));
  assign new_n4303_ = ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & new_n2967_ & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign new_n4304_ = (~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN)) & (P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN) & (~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | (P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN));
  assign new_n4305_ = new_n3191_ & ((P2_STATE2_REG_2__SCAN_IN & (new_n1843_ | new_n4303_)) | ((new_n4301_ | ~P2_STATEBS16_REG_SCAN_IN) & new_n4304_ & ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN));
  assign new_n4306_ = (~new_n4146_ | ~new_n3193_) & (~new_n4303_ | new_n1317_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n4307_ = (new_n2998_ | (new_n4213_ & new_n2996_)) & ~new_n3506_ & ~new_n3353_ & (~new_n2985_ | ~new_n2990_ | new_n2133_);
  assign new_n4308_ = (new_n4309_ | ~new_n4310_ | (~new_n4300_ & P2_INSTQUEUE_REG_4__2__SCAN_IN)) & (new_n4313_ | ~new_n4314_ | (~new_n4300_ & P2_INSTQUEUE_REG_4__4__SCAN_IN));
  assign new_n4309_ = new_n3114_ & ((P2_STATE2_REG_2__SCAN_IN & (new_n1843_ | new_n4303_)) | ((new_n4301_ | ~P2_STATEBS16_REG_SCAN_IN) & new_n4304_ & ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN));
  assign new_n4310_ = new_n4311_ & (~new_n3393_ | ~new_n3189_);
  assign new_n4311_ = ~new_n4312_ & (~new_n3188_ | ~new_n3059_ | (new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) | (~new_n1412_ ^ (new_n1409_ ^ ~new_n1421_)));
  assign new_n4312_ = new_n4303_ & ~new_n1367_ & new_n2966_ & P2_STATE2_REG_3__SCAN_IN;
  assign new_n4313_ = new_n3071_ & ((P2_STATE2_REG_2__SCAN_IN & (new_n1843_ | new_n4303_)) | ((new_n4301_ | ~P2_STATEBS16_REG_SCAN_IN) & new_n4304_ & ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN));
  assign new_n4314_ = new_n4315_ & (~new_n3393_ | ~new_n3069_);
  assign new_n4315_ = ~new_n4316_ & (~new_n3070_ | ~new_n3059_ | (new_n1664_ ^ ((~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_)))) | (~new_n1412_ ^ (new_n1409_ ^ ~new_n1421_)));
  assign new_n4316_ = new_n4303_ & ~new_n1350_ & new_n2966_ & P2_STATE2_REG_3__SCAN_IN;
  assign new_n4317_ = ~new_n4318_ & (new_n4319_ | new_n4320_ | ~new_n4321_) & ~new_n4322_ & (new_n4323_ | new_n4324_ | ~new_n4325_);
  assign new_n4318_ = new_n3109_ & ~new_n4250_;
  assign new_n4319_ = P2_INSTQUEUE_REG_4__1__SCAN_IN & (~new_n4302_ | (~new_n4304_ & (new_n2969_ | (new_n4301_ & new_n2968_))));
  assign new_n4320_ = new_n3115_ & ((P2_STATE2_REG_2__SCAN_IN & (new_n1843_ | new_n4303_)) | ((new_n4301_ | ~P2_STATEBS16_REG_SCAN_IN) & new_n4304_ & ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN));
  assign new_n4321_ = (~new_n3393_ | ~new_n3244_) & (~new_n4146_ | ~new_n3241_) & (~new_n4303_ | new_n1322_ | ~new_n2966_ | ~P2_STATE2_REG_3__SCAN_IN);
  assign new_n4322_ = P1_INSTQUEUE_REG_13__7__SCAN_IN & (~new_n4226_ | (new_n4225_ & (new_n2998_ | (~new_n3378_ & new_n2996_))));
  assign new_n4323_ = P2_INSTQUEUE_REG_10__3__SCAN_IN & (~new_n4181_ | ((new_n1418_ | ~new_n3364_) & (new_n2969_ | (~new_n4180_ & new_n2968_))));
  assign new_n4324_ = new_n3166_ & (new_n4280_ | new_n4281_);
  assign new_n4325_ = ~new_n4326_ & (~new_n4269_ | ~new_n3211_) & (~new_n3273_ | ~new_n2968_ | ~new_n3210_);
  assign new_n4326_ = new_n3538_ & ~new_n1345_ & new_n2966_ & P2_STATE2_REG_3__SCAN_IN;
  assign new_n4327_ = new_n4328_ & new_n4332_ & new_n4343_ & ~new_n4341_ & (~new_n4338_ | (~new_n4265_ & P2_INSTQUEUE_REG_9__7__SCAN_IN));
  assign new_n4328_ = (new_n4331_ | (new_n4208_ & (~new_n4206_ | new_n4207_))) & (~new_n4330_ | ((~new_n2282_ | ~new_n4329_) & new_n2504_ & (new_n2282_ | new_n4329_)));
  assign new_n4329_ = (new_n2237_ & (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_))))) ^ (new_n2279_ ? new_n2281_ : ~new_n2275_);
  assign new_n4330_ = (new_n2505_ | ~P1_EAX_REG_3__SCAN_IN) & (~new_n2505_ | new_n2512_ | (new_n2954_ ? ~BUF1_REG_3__SCAN_IN : ~DATAI_3_));
  assign new_n4331_ = ~P1_INSTQUEUE_REG_4__7__SCAN_IN & ~P1_INSTQUEUE_REG_4__1__SCAN_IN;
  assign new_n4332_ = (~new_n3049_ | (~new_n4333_ & (~P1_STATE2_REG_2__SCAN_IN | ~new_n2120_ | P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN))) & (new_n4335_ | (~new_n4336_ & (~new_n2120_ | ~P1_STATE2_REG_2__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN)));
  assign new_n4333_ = new_n4334_ & (~P1_STATEBS16_REG_SCAN_IN | (new_n2994_ ? ((~new_n2277_ & (new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_))) | (new_n2277_ & ((~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_)))) | new_n2284_ | (~new_n2154_ ^ (~new_n2148_ ^ ~new_n2200_))) : (~new_n2284_ | (~new_n2277_ & (new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_))) | (new_n2277_ & ((~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_)))) | (~new_n2154_ ^ (~new_n2148_ ^ ~new_n2200_)))));
  assign new_n4334_ = new_n2576_ & (new_n4235_ | ((new_n2133_ | new_n2131_ | ((new_n2050_ | new_n2143_) & (~new_n2121_ | (new_n2050_ & new_n2143_)))) & (~new_n2133_ | (~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_))))) & (new_n2131_ ^ ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))) & ~new_n2987_ & (new_n2121_ ^ (new_n2050_ ^ new_n2143_))));
  assign new_n4335_ = (~new_n3003_ | (new_n2954_ & ~BUF1_REG_6__SCAN_IN) | (~new_n2954_ & ~DATAI_6_)) & (~new_n3003_ | (new_n2954_ ? ~BUF1_REG_1__SCAN_IN : ~DATAI_1_));
  assign new_n4336_ = new_n4337_ & (~P1_STATEBS16_REG_SCAN_IN | (new_n2994_ ? ((~new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) | new_n2284_ | (~new_n2154_ ^ (~new_n2148_ ^ ~new_n2200_))) : (~new_n2284_ | (~new_n2277_ ^ ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) | (~new_n2154_ ^ (~new_n2148_ ^ ~new_n2200_)))));
  assign new_n4337_ = new_n2576_ & (new_n2991_ | ((new_n2133_ ^ (~new_n2131_ & ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_))))) & (new_n2131_ ^ ((~new_n2050_ & ~new_n2143_) | (new_n2121_ & (~new_n2050_ | ~new_n2143_)))) & ~new_n2987_ & (new_n2121_ ^ (new_n2050_ ^ new_n2143_))));
  assign new_n4338_ = new_n4339_ & (~new_n4270_ | ~new_n4083_) & (~new_n3113_ | (~new_n4271_ & (~new_n4274_ | (P2_STATEBS16_REG_SCAN_IN & (new_n4269_ | new_n4270_)))));
  assign new_n4339_ = ~new_n4340_ & (~new_n2968_ | ~new_n3274_ | ~new_n2963_ | (new_n1664_ & (~new_n1409_ | new_n1421_) & (~new_n1412_ | (~new_n1409_ & new_n1421_))) | (~new_n1664_ & ((new_n1409_ & ~new_n1421_) | (new_n1412_ & (new_n1409_ | ~new_n1421_)))) | (~new_n1412_ ^ (~new_n1409_ ^ new_n1421_)));
  assign new_n4340_ = ~new_n1335_ & new_n2966_ & P2_STATE2_REG_3__SCAN_IN & new_n3364_ & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign new_n4341_ = (P1_INSTQUEUE_REG_0__1__SCAN_IN | P1_INSTQUEUE_REG_0__7__SCAN_IN) & (~new_n4342_ | (new_n4218_ & (new_n2998_ | (new_n2996_ & ~new_n3161_ & ~new_n4098_))));
  assign new_n4342_ = new_n3003_ & (~P1_STATE2_REG_2__SCAN_IN | ((P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)) & (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ^ ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)))) & (~P1_STATE2_REG_3__SCAN_IN | (~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN));
  assign new_n4343_ = (~P1_INSTQUEUE_REG_6__1__SCAN_IN | (new_n4190_ & (~new_n3041_ | new_n4189_))) & (~P1_INSTQUEUE_REG_8__6__SCAN_IN | (new_n4194_ & (~new_n3032_ | new_n4193_)));
  assign new_n4344_ = (new_n4345_ | ~new_n4349_) & (~new_n2678_ | (~new_n1528_ & new_n1626_) | (new_n1528_ & ~new_n1626_));
  assign new_n4345_ = new_n2649_ & (~new_n4348_ | (~new_n4347_ & (new_n4346_ | new_n2952_))) & (new_n4348_ | new_n4347_ | (~new_n4346_ & ~new_n2952_));
  assign new_n4346_ = ~new_n2263_ & (~new_n2261_ | ~new_n2237_);
  assign new_n4347_ = new_n2263_ & new_n2261_ & new_n2237_;
  assign new_n4348_ = ~new_n2258_ ^ (new_n2237_ & (~new_n2257_ | (~new_n2198_ & (new_n2251_ | new_n2185_))) & (new_n2257_ | new_n2198_ | (~new_n2251_ & ~new_n2185_)));
  assign new_n4349_ = (~new_n2639_ | (~new_n2647_ & ~P1_REIP_REG_6__SCAN_IN) | (new_n2647_ & P1_REIP_REG_6__SCAN_IN)) & (~new_n2643_ | ~new_n2259_) & new_n4350_ & (new_n2640_ | ~P1_EBX_REG_6__SCAN_IN);
  assign new_n4350_ = (~new_n2629_ | ~new_n2769_) & ~new_n2636_ & (~new_n2630_ | ~P1_REIP_REG_6__SCAN_IN) & (~P1_PHYADDRPOINTER_REG_6__SCAN_IN | new_n2630_ | ~P1_STATE2_REG_3__SCAN_IN);
  assign new_n4351_ = ~new_n4352_ & ((new_n1646_ & new_n2683_ & ~new_n1335_) | (~new_n2683_ & P2_EBX_REG_19__SCAN_IN) | ((new_n2765_ | ~new_n1997_) & new_n2683_ & new_n1335_ & (~new_n2765_ | new_n1997_)));
  assign new_n4352_ = new_n4353_ & ((~new_n1655_ & ~new_n1683_ & (new_n1684_ | (~new_n1651_ ^ ~new_n1428_)) & (~new_n1684_ | (~new_n1651_ & ~new_n1428_) | (new_n1651_ & new_n1428_))) | ~new_n1758_ | ((new_n1655_ | new_n1683_) & (new_n1684_ ^ (new_n1651_ ^ ~new_n1428_))));
  assign new_n4353_ = (~new_n1684_ | ~new_n1759_ | ~new_n1335_) & (new_n1759_ | ~P2_EAX_REG_11__SCAN_IN) & (new_n1784_ | ~new_n1759_ | new_n1335_ | (~new_n2976_ & ~BUF2_REG_11__SCAN_IN) | (new_n2976_ & ~BUF1_REG_11__SCAN_IN));
  assign new_n4354_ = new_n4355_ & ~new_n4400_ & ((new_n4397_ & new_n2040_) | new_n4399_ | ~new_n4413_ | (new_n2004_ & new_n3313_));
  assign new_n4355_ = new_n4358_ & ((~new_n4356_ & ~new_n4357_) | ~new_n1758_ | (new_n4356_ & new_n4357_)) & new_n4388_ & ~new_n4359_ & new_n4360_ & new_n4382_;
  assign new_n4356_ = (new_n1658_ | new_n1681_) & ((new_n1658_ & new_n1681_) | (~new_n1659_ & (~new_n1680_ | (new_n1677_ & (new_n1661_ | ~new_n1675_)))));
  assign new_n4357_ = ~new_n1656_ & ~new_n1683_;
  assign new_n4358_ = (~new_n2678_ | (~new_n1529_ & new_n1625_) | (new_n1529_ & ~new_n1625_)) & (~new_n2690_ | (~new_n2002_ & ~new_n2001_ & new_n1976_ & ~new_n2000_) | (new_n2002_ & (new_n2001_ | ~new_n1976_ | new_n2000_)));
  assign new_n4359_ = new_n2604_ & ((~new_n2533_ & P1_INSTADDRPOINTER_REG_6__SCAN_IN) | (new_n2533_ & ~P1_INSTADDRPOINTER_REG_6__SCAN_IN) | ((new_n2534_ | ~P1_INSTADDRPOINTER_REG_5__SCAN_IN) & (new_n2535_ | (new_n2534_ & ~P1_INSTADDRPOINTER_REG_5__SCAN_IN)))) & ((~new_n2533_ ^ P1_INSTADDRPOINTER_REG_6__SCAN_IN) | (~new_n2534_ & P1_INSTADDRPOINTER_REG_5__SCAN_IN) | (~new_n2535_ & (~new_n2534_ | P1_INSTADDRPOINTER_REG_5__SCAN_IN)));
  assign new_n4360_ = ~new_n4361_ & ~new_n4381_ & (new_n4366_ | ~new_n4371_) & ~new_n4376_ & (new_n4377_ | ~new_n4378_);
  assign new_n4361_ = (new_n4362_ | ~new_n2937_) & (~P3_INSTADDRPOINTER_REG_24__SCAN_IN | new_n2937_ | new_n3282_) & (~P3_REIP_REG_24__SCAN_IN | P3_STATE2_REG_2__SCAN_IN | (~new_n2937_ & ~new_n3282_));
  assign new_n4362_ = new_n4363_ & (((~new_n2925_ ^ ~P3_INSTADDRPOINTER_REG_24__SCAN_IN) & ((new_n2925_ & ~P3_INSTADDRPOINTER_REG_23__SCAN_IN) | ~new_n2930_ | (new_n2925_ & ~P3_INSTADDRPOINTER_REG_22__SCAN_IN)) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_23__SCAN_IN) & (new_n2925_ | new_n2936_) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN)) | ~new_n2935_ | ((~new_n2925_ | P3_INSTADDRPOINTER_REG_24__SCAN_IN) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_24__SCAN_IN) & (((~new_n2925_ | P3_INSTADDRPOINTER_REG_23__SCAN_IN) & new_n2930_ & (~new_n2925_ | P3_INSTADDRPOINTER_REG_22__SCAN_IN)) | (~new_n2925_ & P3_INSTADDRPOINTER_REG_23__SCAN_IN) | (~new_n2925_ & ~new_n2936_) | (~new_n2925_ & P3_INSTADDRPOINTER_REG_22__SCAN_IN))));
  assign new_n4363_ = ((~P3_INSTADDRPOINTER_REG_24__SCAN_IN & (~P3_INSTADDRPOINTER_REG_23__SCAN_IN | ~new_n2864_ | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN)) | ~new_n2928_ | (P3_INSTADDRPOINTER_REG_24__SCAN_IN & P3_INSTADDRPOINTER_REG_23__SCAN_IN & new_n2864_ & P3_INSTADDRPOINTER_REG_22__SCAN_IN)) & new_n4364_ & ((~P3_INSTADDRPOINTER_REG_24__SCAN_IN & (~P3_INSTADDRPOINTER_REG_23__SCAN_IN | ~new_n2912_ | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN)) | ~new_n2926_ | (P3_INSTADDRPOINTER_REG_24__SCAN_IN & P3_INSTADDRPOINTER_REG_23__SCAN_IN & new_n2912_ & P3_INSTADDRPOINTER_REG_22__SCAN_IN));
  assign new_n4364_ = new_n4365_ & (new_n4205_ | (new_n2851_ & P3_INSTADDRPOINTER_REG_0__SCAN_IN) | (~P3_INSTADDRPOINTER_REG_24__SCAN_IN & (~new_n2842_ | ~P3_INSTADDRPOINTER_REG_23__SCAN_IN)));
  assign new_n4365_ = (new_n3287_ | (~P3_INSTADDRPOINTER_REG_24__SCAN_IN & (~P3_INSTADDRPOINTER_REG_23__SCAN_IN | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN | ~new_n2780_ | ~new_n2786_)) | (P3_INSTADDRPOINTER_REG_24__SCAN_IN & P3_INSTADDRPOINTER_REG_23__SCAN_IN & P3_INSTADDRPOINTER_REG_22__SCAN_IN & new_n2780_ & new_n2786_)) & (~new_n2850_ | (P3_INSTADDRPOINTER_REG_24__SCAN_IN & P3_INSTADDRPOINTER_REG_23__SCAN_IN & P3_INSTADDRPOINTER_REG_22__SCAN_IN & new_n2848_ & new_n2786_) | (~P3_INSTADDRPOINTER_REG_24__SCAN_IN & (~P3_INSTADDRPOINTER_REG_23__SCAN_IN | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN | ~new_n2848_ | ~new_n2786_)));
  assign new_n4366_ = P1_INSTQUEUE_REG_12__5__SCAN_IN & (~new_n4370_ | (new_n4368_ & (new_n2998_ | (new_n2996_ & ~new_n3120_ & ~new_n4367_))));
  assign new_n4367_ = new_n2284_ & new_n2994_ & (new_n2277_ | (~new_n2148_ & ~new_n2200_) | (~new_n2154_ & (~new_n2148_ | ~new_n2200_))) & (~new_n2277_ | ((new_n2148_ | new_n2200_) & (new_n2154_ | (new_n2148_ & new_n2200_)))) & (new_n2154_ ^ (new_n2148_ ^ new_n2200_));
  assign new_n4368_ = ~new_n4369_ & (~new_n2986_ | new_n2987_ | ~new_n2990_ | new_n2133_);
  assign new_n4369_ = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign new_n4370_ = new_n3003_ & (~P1_STATE2_REG_2__SCAN_IN | (P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ^ ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)))) & (~P1_STATE2_REG_3__SCAN_IN | (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN));
  assign new_n4371_ = (~new_n3053_ | (~new_n4375_ & (~new_n4372_ | (P1_STATEBS16_REG_SCAN_IN & (new_n3120_ | new_n4367_))))) & new_n4373_ & (~new_n4367_ | ~new_n3054_);
  assign new_n4372_ = new_n2576_ & (new_n4369_ | (new_n2986_ & ~new_n2987_ & new_n2990_ & ~new_n2133_));
  assign new_n4373_ = ~new_n4374_ & (~new_n3055_ | new_n2994_ | (~new_n2277_ & (new_n2154_ | (new_n2148_ & new_n2200_)) & (new_n2148_ | new_n2200_)) | (new_n2277_ & ((~new_n2154_ & (~new_n2148_ | ~new_n2200_)) | (~new_n2148_ & ~new_n2200_))) | new_n2284_ | (~new_n2154_ & (~new_n2148_ | ~new_n2200_) & (new_n2148_ | new_n2200_)) | (new_n2154_ & (~new_n2148_ ^ new_n2200_)));
  assign new_n4374_ = new_n3056_ & new_n4369_;
  assign new_n4375_ = P1_STATE2_REG_2__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & (~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ^ P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN) & (P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | (P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN)) & (~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  assign new_n4376_ = (~new_n1998_ | (~new_n1997_ & ~new_n1996_ & ~new_n1995_ & ~new_n1994_ & new_n1977_ & ~new_n1993_)) & new_n2691_ & (new_n1998_ | new_n1997_ | new_n1996_ | new_n1995_ | new_n1994_ | ~new_n1977_ | new_n1993_);
  assign new_n4377_ = P1_INSTQUEUE_REG_12__6__SCAN_IN & (~new_n4370_ | (new_n4368_ & (new_n2998_ | (new_n2996_ & ~new_n3120_ & ~new_n4367_))));
  assign new_n4378_ = (~new_n3048_ | (~new_n4375_ & (~new_n4372_ | (P1_STATEBS16_REG_SCAN_IN & (new_n3120_ | new_n4367_))))) & new_n4379_ & (~new_n4367_ | ~new_n3165_);
  assign new_n4379_ = ~new_n4380_ & (~new_n3119_ | new_n2994_ | (~new_n2277_ & (new_n2154_ | (new_n2148_ & new_n2200_)) & (new_n2148_ | new_n2200_)) | (new_n2277_ & ((~new_n2154_ & (~new_n2148_ | ~new_n2200_)) | (~new_n2148_ & ~new_n2200_))) | new_n2284_ | (~new_n2154_ & (~new_n2148_ | ~new_n2200_) & (new_n2148_ | new_n2200_)) | (new_n2154_ & (~new_n2148_ ^ new_n2200_)));
  assign new_n4380_ = new_n3351_ & new_n4369_;
  assign new_n4381_ = ((~new_n2925_ & ~P3_INSTADDRPOINTER_REG_21__SCAN_IN) | (new_n2925_ & P3_INSTADDRPOINTER_REG_21__SCAN_IN) | (~new_n2925_ & (~new_n4241_ | P3_INSTADDRPOINTER_REG_19__SCAN_IN)) | (P3_INSTADDRPOINTER_REG_20__SCAN_IN & (~new_n2925_ | (~new_n4241_ & P3_INSTADDRPOINTER_REG_19__SCAN_IN)))) & new_n3289_ & ((~new_n2925_ ^ ~P3_INSTADDRPOINTER_REG_21__SCAN_IN) | ((new_n2925_ | (new_n4241_ & ~P3_INSTADDRPOINTER_REG_19__SCAN_IN)) & (~P3_INSTADDRPOINTER_REG_20__SCAN_IN | (new_n2925_ & (new_n4241_ | ~P3_INSTADDRPOINTER_REG_19__SCAN_IN)))));
  assign new_n4382_ = (~new_n4383_ | (new_n1694_ & new_n2665_)) & ((~new_n1976_ & new_n2000_) | ~new_n2691_ | (new_n1976_ & ~new_n2000_));
  assign new_n4383_ = new_n4384_ & ((new_n1996_ & (new_n1995_ | new_n1994_ | ~new_n1977_ | new_n1993_)) | ~new_n2691_ | (~new_n1996_ & ~new_n1995_ & ~new_n1994_ & new_n1977_ & ~new_n1993_));
  assign new_n4384_ = ~new_n4385_ & ~new_n4386_ & (~new_n2757_ | (~new_n1939_ & ~new_n1940_) | (new_n1939_ & new_n1940_)) & new_n4387_ & (new_n2723_ | ~P2_EBX_REG_18__SCAN_IN);
  assign new_n4385_ = ~new_n2727_ & ~new_n2724_ & P2_STATE2_REG_1__SCAN_IN & (~new_n2735_ | ~new_n2736_ | ~new_n2751_) & (new_n2735_ | (new_n2736_ & new_n2751_));
  assign new_n4386_ = (new_n2732_ | P2_PHYADDRPOINTER_REG_18__SCAN_IN) & (~new_n2732_ | ~P2_PHYADDRPOINTER_REG_18__SCAN_IN) & new_n2727_ & ~new_n2724_ & P2_STATE2_REG_1__SCAN_IN;
  assign new_n4387_ = (~P2_PHYADDRPOINTER_REG_18__SCAN_IN | new_n2724_ | ~P2_STATE2_REG_3__SCAN_IN) & (~new_n2724_ | ~P2_REIP_REG_18__SCAN_IN) & (new_n2724_ | ~new_n3374_);
  assign new_n4388_ = ~new_n4389_ & (~new_n2602_ | (new_n4348_ & (new_n4347_ | (~new_n4346_ & ~new_n2952_))) | (~new_n4348_ & ~new_n4347_ & (new_n4346_ | new_n2952_)));
  assign new_n4389_ = new_n4396_ & (~new_n2937_ | (new_n4391_ & (((~new_n4390_ | (~new_n2925_ & P3_INSTADDRPOINTER_REG_25__SCAN_IN)) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_26__SCAN_IN) & (~new_n2925_ | (P3_INSTADDRPOINTER_REG_25__SCAN_IN & P3_INSTADDRPOINTER_REG_26__SCAN_IN))) | ~new_n2935_ | ((new_n4390_ | (new_n2925_ & ~P3_INSTADDRPOINTER_REG_25__SCAN_IN)) & (~P3_INSTADDRPOINTER_REG_25__SCAN_IN | ~P3_INSTADDRPOINTER_REG_26__SCAN_IN) & (new_n2925_ ^ P3_INSTADDRPOINTER_REG_26__SCAN_IN)))));
  assign new_n4390_ = ((new_n2925_ & ~P3_INSTADDRPOINTER_REG_24__SCAN_IN) | (new_n2925_ & ~P3_INSTADDRPOINTER_REG_23__SCAN_IN) | ~new_n2930_ | (new_n2925_ & ~P3_INSTADDRPOINTER_REG_22__SCAN_IN)) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_24__SCAN_IN) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_23__SCAN_IN) & (new_n2925_ | new_n2936_) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  assign new_n4391_ = ~new_n4392_ & ~new_n4393_ & new_n4394_ & (new_n4395_ | (~P3_INSTADDRPOINTER_REG_26__SCAN_IN & (~P3_INSTADDRPOINTER_REG_25__SCAN_IN | ~new_n2851_ | ~P3_INSTADDRPOINTER_REG_0__SCAN_IN)) | (P3_INSTADDRPOINTER_REG_26__SCAN_IN & P3_INSTADDRPOINTER_REG_25__SCAN_IN & new_n2851_ & P3_INSTADDRPOINTER_REG_0__SCAN_IN));
  assign new_n4392_ = (P3_INSTADDRPOINTER_REG_26__SCAN_IN | (P3_INSTADDRPOINTER_REG_25__SCAN_IN & P3_INSTADDRPOINTER_REG_24__SCAN_IN & P3_INSTADDRPOINTER_REG_23__SCAN_IN & new_n2864_ & P3_INSTADDRPOINTER_REG_22__SCAN_IN)) & new_n2928_ & (~P3_INSTADDRPOINTER_REG_25__SCAN_IN | ~P3_INSTADDRPOINTER_REG_26__SCAN_IN | ~P3_INSTADDRPOINTER_REG_24__SCAN_IN | ~P3_INSTADDRPOINTER_REG_23__SCAN_IN | ~new_n2864_ | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  assign new_n4393_ = (P3_INSTADDRPOINTER_REG_26__SCAN_IN | (P3_INSTADDRPOINTER_REG_25__SCAN_IN & P3_INSTADDRPOINTER_REG_24__SCAN_IN & P3_INSTADDRPOINTER_REG_23__SCAN_IN & new_n2912_ & P3_INSTADDRPOINTER_REG_22__SCAN_IN)) & new_n2926_ & (~P3_INSTADDRPOINTER_REG_25__SCAN_IN | ~P3_INSTADDRPOINTER_REG_26__SCAN_IN | ~P3_INSTADDRPOINTER_REG_24__SCAN_IN | ~P3_INSTADDRPOINTER_REG_23__SCAN_IN | ~new_n2912_ | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  assign new_n4394_ = (new_n3287_ | (P3_INSTADDRPOINTER_REG_26__SCAN_IN & new_n2851_ & P3_INSTADDRPOINTER_REG_25__SCAN_IN) | (~P3_INSTADDRPOINTER_REG_26__SCAN_IN & (~new_n2851_ | ~P3_INSTADDRPOINTER_REG_25__SCAN_IN))) & (~new_n2850_ | (~P3_INSTADDRPOINTER_REG_26__SCAN_IN & (~new_n2847_ | ~P3_INSTADDRPOINTER_REG_25__SCAN_IN)) | (new_n2847_ & P3_INSTADDRPOINTER_REG_25__SCAN_IN & P3_INSTADDRPOINTER_REG_26__SCAN_IN)) & ((P3_INSTADDRPOINTER_REG_26__SCAN_IN & P3_INSTADDRPOINTER_REG_25__SCAN_IN & new_n2851_ & P3_INSTADDRPOINTER_REG_0__SCAN_IN) | ~new_n2845_ | (~P3_INSTADDRPOINTER_REG_26__SCAN_IN & (~P3_INSTADDRPOINTER_REG_25__SCAN_IN | ~new_n2851_ | ~P3_INSTADDRPOINTER_REG_0__SCAN_IN)));
  assign new_n4395_ = (new_n2809_ | ~new_n2802_ | ~new_n2790_ | ~new_n2821_ | ~new_n2826_ | ~new_n2833_ | ~new_n2796_ | new_n2815_) & (new_n2802_ | ~new_n2809_ | ~new_n2833_ | new_n2790_ | new_n2796_ | ~new_n2815_ | new_n2826_ | new_n2821_) & (~new_n2826_ | ~new_n2821_ | ~new_n2833_ | new_n2790_ | new_n2796_ | new_n2815_ | new_n2802_ | ~new_n2809_) & (~new_n2790_ | ~new_n2821_ | ~new_n2802_ | ~new_n2809_ | new_n2826_ | ~new_n2815_ | new_n2833_) & (~new_n2815_ | ((~new_n2802_ | new_n2809_ | (~new_n2821_ & (~new_n2790_ | new_n2796_) & ~new_n2826_ & (new_n2790_ | ~new_n2796_))) & (~new_n2809_ | ((~new_n2790_ | ~new_n2833_) & (~new_n2802_ | new_n2790_ | new_n2796_))) & ((new_n2796_ & new_n2826_) | new_n2802_ | (~new_n2826_ & ~new_n2821_)))) & (new_n2796_ | ~new_n2821_ | (new_n2809_ & (~new_n2802_ | ~new_n2826_))) & (new_n2796_ | new_n2802_ | ~new_n2790_ | ~new_n2833_) & (new_n2802_ | ~new_n2790_ | ~new_n2826_) & ((~new_n2790_ & ~new_n2796_) | new_n2802_ | ~new_n2809_) & (~new_n2796_ | new_n2821_ | (new_n2790_ & new_n2833_)) & (new_n2833_ | ((~new_n2802_ | new_n2809_) & ~new_n2826_ & (new_n2790_ | new_n2796_))) & (new_n2815_ | (new_n2821_ & (new_n2790_ ? new_n2826_ : ~new_n2796_))) & ((new_n2802_ ^ new_n2809_) | ~new_n2826_ | ~new_n2833_ | ~new_n2815_ | ~new_n2821_ | new_n2790_ | ~new_n2796_);
  assign new_n4396_ = (~new_n3997_ | ~P3_INSTADDRPOINTER_REG_26__SCAN_IN) & (~P3_REIP_REG_26__SCAN_IN | new_n3997_ | P3_STATE2_REG_2__SCAN_IN);
  assign new_n4397_ = new_n4398_ ^ ((~new_n1890_ & P2_INSTADDRPOINTER_REG_4__SCAN_IN) | ((~new_n1903_ | (~new_n1892_ & P2_INSTADDRPOINTER_REG_3__SCAN_IN)) & (~new_n1892_ | P2_INSTADDRPOINTER_REG_3__SCAN_IN) & (~new_n1890_ | P2_INSTADDRPOINTER_REG_4__SCAN_IN)));
  assign new_n4398_ = P2_INSTADDRPOINTER_REG_5__SCAN_IN ^ (new_n1887_ | (new_n1534_ & (new_n1860_ | new_n1855_ | ~new_n1820_ | ~new_n1849_) & (~new_n1860_ | (~new_n1855_ & new_n1820_ & new_n1849_))));
  assign new_n4399_ = new_n2028_ & ((new_n1962_ & P2_INSTADDRPOINTER_REG_5__SCAN_IN) | (~new_n1962_ & ~P2_INSTADDRPOINTER_REG_5__SCAN_IN) | ((~new_n1963_ | ~P2_INSTADDRPOINTER_REG_4__SCAN_IN) & ((~new_n1963_ & ~P2_INSTADDRPOINTER_REG_4__SCAN_IN) | ((~new_n1964_ | ~P2_INSTADDRPOINTER_REG_3__SCAN_IN) & (~new_n1965_ | (~new_n1964_ & ~P2_INSTADDRPOINTER_REG_3__SCAN_IN)))))) & ((new_n1962_ ^ P2_INSTADDRPOINTER_REG_5__SCAN_IN) | (new_n1963_ & P2_INSTADDRPOINTER_REG_4__SCAN_IN) | ((new_n1963_ | P2_INSTADDRPOINTER_REG_4__SCAN_IN) & ((new_n1964_ & P2_INSTADDRPOINTER_REG_3__SCAN_IN) | (new_n1965_ & (new_n1964_ | P2_INSTADDRPOINTER_REG_3__SCAN_IN)))));
  assign new_n4400_ = new_n2937_ & (new_n4401_ | ~new_n4403_);
  assign new_n4401_ = (P3_INSTADDRPOINTER_REG_31__SCAN_IN | (((~new_n4402_ & new_n2923_ & P3_INSTADDRPOINTER_REG_29__SCAN_IN & P3_INSTADDRPOINTER_REG_27__SCAN_IN & P3_INSTADDRPOINTER_REG_28__SCAN_IN) | P3_INSTADDRPOINTER_REG_30__SCAN_IN | (~new_n2923_ & ~P3_INSTADDRPOINTER_REG_29__SCAN_IN & ~P3_INSTADDRPOINTER_REG_27__SCAN_IN & ~P3_INSTADDRPOINTER_REG_28__SCAN_IN)) & (~new_n4402_ | ~P3_INSTADDRPOINTER_REG_30__SCAN_IN | new_n2923_ | P3_INSTADDRPOINTER_REG_29__SCAN_IN | P3_INSTADDRPOINTER_REG_27__SCAN_IN | P3_INSTADDRPOINTER_REG_28__SCAN_IN))) & new_n2935_ & (new_n4402_ | (new_n2923_ ? (~P3_INSTADDRPOINTER_REG_30__SCAN_IN | ~P3_INSTADDRPOINTER_REG_31__SCAN_IN | ~P3_INSTADDRPOINTER_REG_29__SCAN_IN | ~P3_INSTADDRPOINTER_REG_27__SCAN_IN | ~P3_INSTADDRPOINTER_REG_28__SCAN_IN) : (P3_INSTADDRPOINTER_REG_30__SCAN_IN | P3_INSTADDRPOINTER_REG_31__SCAN_IN)));
  assign new_n4402_ = (new_n2925_ | ~P3_INSTADDRPOINTER_REG_25__SCAN_IN) & (new_n2925_ | ~P3_INSTADDRPOINTER_REG_26__SCAN_IN) & (new_n4390_ | (new_n2925_ & (~P3_INSTADDRPOINTER_REG_25__SCAN_IN | ~P3_INSTADDRPOINTER_REG_26__SCAN_IN)));
  assign new_n4403_ = ((P3_INSTADDRPOINTER_REG_31__SCAN_IN & new_n4404_ & P3_INSTADDRPOINTER_REG_30__SCAN_IN) | ~new_n2928_ | (~P3_INSTADDRPOINTER_REG_31__SCAN_IN & (~new_n4404_ | ~P3_INSTADDRPOINTER_REG_30__SCAN_IN))) & ((~new_n4404_ & ~P3_INSTADDRPOINTER_REG_30__SCAN_IN) | ~new_n2928_ | (new_n4404_ & P3_INSTADDRPOINTER_REG_30__SCAN_IN)) & new_n4407_ & ~new_n4412_ & ((~new_n4406_ & ~P3_INSTADDRPOINTER_REG_30__SCAN_IN & ~P3_INSTADDRPOINTER_REG_31__SCAN_IN) | ~new_n2926_ | (new_n4406_ & P3_INSTADDRPOINTER_REG_30__SCAN_IN & P3_INSTADDRPOINTER_REG_31__SCAN_IN));
  assign new_n4404_ = new_n4405_ & P3_INSTADDRPOINTER_REG_26__SCAN_IN & P3_INSTADDRPOINTER_REG_25__SCAN_IN & P3_INSTADDRPOINTER_REG_24__SCAN_IN & new_n2863_ & P3_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign new_n4405_ = P3_INSTADDRPOINTER_REG_29__SCAN_IN & P3_INSTADDRPOINTER_REG_27__SCAN_IN & P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign new_n4406_ = new_n4405_ & P3_INSTADDRPOINTER_REG_26__SCAN_IN & P3_INSTADDRPOINTER_REG_25__SCAN_IN & P3_INSTADDRPOINTER_REG_24__SCAN_IN & new_n2911_ & P3_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign new_n4407_ = new_n4408_ & ((P3_INSTADDRPOINTER_REG_30__SCAN_IN & P3_INSTADDRPOINTER_REG_31__SCAN_IN & new_n4411_ & new_n4405_) | ~new_n2845_ | ((~new_n4411_ | ~new_n4405_) & ~P3_INSTADDRPOINTER_REG_30__SCAN_IN & ~P3_INSTADDRPOINTER_REG_31__SCAN_IN));
  assign new_n4408_ = (new_n4410_ | ~new_n2850_) & ((P3_INSTADDRPOINTER_REG_31__SCAN_IN & new_n4409_ & new_n4405_ & P3_INSTADDRPOINTER_REG_30__SCAN_IN) | new_n3553_ | (~P3_INSTADDRPOINTER_REG_31__SCAN_IN & (~new_n4409_ | ~new_n4405_ | ~P3_INSTADDRPOINTER_REG_30__SCAN_IN))) & (new_n3287_ | (~P3_INSTADDRPOINTER_REG_30__SCAN_IN & (~new_n4409_ | ~new_n4405_)) | (new_n4409_ & new_n4405_ & P3_INSTADDRPOINTER_REG_30__SCAN_IN));
  assign new_n4409_ = P3_INSTADDRPOINTER_REG_26__SCAN_IN & new_n2851_ & P3_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign new_n4410_ = (P3_INSTADDRPOINTER_REG_31__SCAN_IN | ((~new_n2847_ | ~P3_INSTADDRPOINTER_REG_25__SCAN_IN | ~new_n4405_ | ~P3_INSTADDRPOINTER_REG_26__SCAN_IN) & (~new_n4405_ | ~P3_INSTADDRPOINTER_REG_30__SCAN_IN | ~new_n2847_ | ~P3_INSTADDRPOINTER_REG_25__SCAN_IN | ~P3_INSTADDRPOINTER_REG_26__SCAN_IN))) & ((~P3_INSTADDRPOINTER_REG_30__SCAN_IN & ~P3_INSTADDRPOINTER_REG_31__SCAN_IN) | (new_n4405_ & P3_INSTADDRPOINTER_REG_30__SCAN_IN & new_n2847_ & P3_INSTADDRPOINTER_REG_25__SCAN_IN & P3_INSTADDRPOINTER_REG_26__SCAN_IN));
  assign new_n4411_ = P3_INSTADDRPOINTER_REG_26__SCAN_IN & P3_INSTADDRPOINTER_REG_25__SCAN_IN & new_n2851_ & P3_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign new_n4412_ = ~new_n4395_ & (~P3_INSTADDRPOINTER_REG_0__SCAN_IN | ~P3_INSTADDRPOINTER_REG_31__SCAN_IN | ~new_n4409_ | ~new_n4405_ | ~P3_INSTADDRPOINTER_REG_30__SCAN_IN) & (P3_INSTADDRPOINTER_REG_30__SCAN_IN | P3_INSTADDRPOINTER_REG_31__SCAN_IN | (P3_INSTADDRPOINTER_REG_0__SCAN_IN & new_n4409_ & new_n4405_));
  assign new_n4413_ = (~P2_REIP_REG_5__SCAN_IN | new_n2005_ | ~new_n2022_) & (~new_n2005_ | ~P2_PHYADDRPOINTER_REG_5__SCAN_IN) & (new_n2005_ | new_n2021_ | (~new_n2743_ & ~P2_PHYADDRPOINTER_REG_5__SCAN_IN) | (new_n2743_ & P2_PHYADDRPOINTER_REG_5__SCAN_IN));
  assign new_n4414_ = ~new_n4415_ & (~new_n4420_ | ((new_n1881_ | new_n1884_ | new_n1798_ | new_n1880_) & new_n4417_ & ((~new_n1881_ & ~new_n1884_) | (~new_n1798_ & ~new_n1880_))));
  assign new_n4415_ = (~new_n4416_ | ((~new_n1650_ | ~new_n1686_) & ((~new_n1650_ & ~new_n1686_) | new_n1652_ | (new_n1685_ & (new_n1655_ | ~new_n1682_))))) & new_n1758_ & (new_n4416_ | (new_n1650_ & new_n1686_) | ((new_n1650_ | new_n1686_) & ~new_n1652_ & (~new_n1685_ | (~new_n1655_ & new_n1682_))));
  assign new_n4416_ = new_n1689_ ^ (new_n1311_ ? new_n1471_ : (new_n1315_ & ~new_n1471_));
  assign new_n4417_ = (~new_n4398_ ^ ((~new_n1890_ & P2_INSTADDRPOINTER_REG_4__SCAN_IN) | ((~new_n1903_ | (P2_INSTADDRPOINTER_REG_3__SCAN_IN & ((~new_n4418_ & P2_INSTADDRPOINTER_REG_2__SCAN_IN) | (new_n4419_ & (~new_n4418_ | P2_INSTADDRPOINTER_REG_2__SCAN_IN))))) & (~new_n1890_ | P2_INSTADDRPOINTER_REG_4__SCAN_IN) & (P2_INSTADDRPOINTER_REG_3__SCAN_IN | (~new_n4418_ & P2_INSTADDRPOINTER_REG_2__SCAN_IN) | (new_n4419_ & (~new_n4418_ | P2_INSTADDRPOINTER_REG_2__SCAN_IN)))))) & (~new_n4419_ | (~new_n4418_ ^ P2_INSTADDRPOINTER_REG_2__SCAN_IN)) & (new_n4419_ | (~new_n4418_ & P2_INSTADDRPOINTER_REG_2__SCAN_IN) | (new_n4418_ & ~P2_INSTADDRPOINTER_REG_2__SCAN_IN));
  assign new_n4418_ = new_n1534_ ? ~new_n1893_ : ~new_n1902_;
  assign new_n4419_ = (new_n1894_ | P2_INSTADDRPOINTER_REG_1__SCAN_IN) & (new_n1900_ | (new_n1894_ & P2_INSTADDRPOINTER_REG_1__SCAN_IN));
  assign new_n4420_ = new_n2705_ & new_n1764_;
  assign new_n4421_ = ((new_n2530_ & (~new_n2525_ ^ ~P1_INSTADDRPOINTER_REG_8__SCAN_IN)) | ~new_n2596_ | (~new_n2530_ & (~new_n2525_ | P1_INSTADDRPOINTER_REG_8__SCAN_IN) & (new_n2525_ | ~P1_INSTADDRPOINTER_REG_8__SCAN_IN))) & new_n4422_ & (~P1_INSTADDRPOINTER_REG_8__SCAN_IN | (~new_n2574_ & (~new_n2588_ | new_n2594_)));
  assign new_n4422_ = (~new_n2589_ | ~P1_REIP_REG_8__SCAN_IN) & new_n4423_ & (~new_n2564_ | ~new_n4424_) & (~new_n2588_ | ~new_n2594_ | P1_INSTADDRPOINTER_REG_8__SCAN_IN);
  assign new_n4423_ = (~new_n2584_ | (~new_n2581_ ^ P1_INSTADDRPOINTER_REG_8__SCAN_IN)) & (~new_n2586_ | (~P1_INSTADDRPOINTER_REG_8__SCAN_IN & ~P1_INSTADDRPOINTER_REG_0__SCAN_IN) | (P1_INSTADDRPOINTER_REG_0__SCAN_IN & (new_n2581_ | ~P1_INSTADDRPOINTER_REG_8__SCAN_IN) & (~new_n2581_ | P1_INSTADDRPOINTER_REG_8__SCAN_IN)));
  assign new_n4424_ = new_n2457_ ^ (~new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_8__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_8__SCAN_IN)));
  assign new_n4425_ = (new_n4427_ | ~new_n4429_ | ((new_n4426_ | ~new_n4428_) & new_n2040_ & (~new_n4426_ | new_n4428_))) & ((new_n1959_ & P2_INSTADDRPOINTER_REG_13__SCAN_IN) | ~new_n2028_ | (~new_n1959_ & ~P2_INSTADDRPOINTER_REG_13__SCAN_IN));
  assign new_n4426_ = ~new_n1798_ & (new_n1880_ | (~new_n1881_ & ~new_n1884_));
  assign new_n4427_ = (((P2_INSTADDRPOINTER_REG_7__SCAN_IN | (~new_n1800_ ^ (new_n1882_ & ~new_n1865_))) & ((P2_INSTADDRPOINTER_REG_7__SCAN_IN & (new_n1800_ | ~new_n1882_ | new_n1865_) & (~new_n1800_ | (new_n1882_ & ~new_n1865_))) | ((P2_INSTADDRPOINTER_REG_6__SCAN_IN | (new_n1882_ ^ ~new_n1865_)) & (new_n1961_ | (P2_INSTADDRPOINTER_REG_6__SCAN_IN & (~new_n1882_ | new_n1865_) & (new_n1882_ | ~new_n1865_)))))) | (~P2_INSTADDRPOINTER_REG_8__SCAN_IN ^ (new_n1800_ | ~new_n1882_ | new_n1865_))) & new_n2028_ & ((~P2_INSTADDRPOINTER_REG_7__SCAN_IN & (new_n1800_ ^ (new_n1882_ & ~new_n1865_))) | ((~P2_INSTADDRPOINTER_REG_7__SCAN_IN | (~new_n1800_ & new_n1882_ & ~new_n1865_) | (new_n1800_ & (~new_n1882_ | new_n1865_))) & ((~P2_INSTADDRPOINTER_REG_6__SCAN_IN & (~new_n1882_ ^ ~new_n1865_)) | (~new_n1961_ & (~P2_INSTADDRPOINTER_REG_6__SCAN_IN | (new_n1882_ & ~new_n1865_) | (~new_n1882_ & new_n1865_))))) | (~P2_INSTADDRPOINTER_REG_8__SCAN_IN & (new_n1800_ | ~new_n1882_ | new_n1865_)) | (P2_INSTADDRPOINTER_REG_8__SCAN_IN & ~new_n1800_ & new_n1882_ & ~new_n1865_));
  assign new_n4428_ = ~P2_INSTADDRPOINTER_REG_8__SCAN_IN ^ (new_n1534_ ? ~new_n1905_ : ~new_n1910_);
  assign new_n4429_ = (~new_n4149_ | ~new_n2004_) & (new_n2005_ | new_n2021_ | (new_n4430_ & P2_PHYADDRPOINTER_REG_8__SCAN_IN) | (~new_n4430_ & ~P2_PHYADDRPOINTER_REG_8__SCAN_IN)) & (~new_n2005_ | ~P2_PHYADDRPOINTER_REG_8__SCAN_IN) & (~P2_REIP_REG_8__SCAN_IN | new_n2005_ | ~new_n2022_);
  assign new_n4430_ = P2_PHYADDRPOINTER_REG_7__SCAN_IN & P2_PHYADDRPOINTER_REG_6__SCAN_IN & new_n2743_ & P2_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign new_n4431_ = ~new_n4432_ & (((new_n1931_ | P2_INSTADDRPOINTER_REG_13__SCAN_IN) & (~new_n1931_ | ~P2_INSTADDRPOINTER_REG_13__SCAN_IN) & ~new_n1797_ & ~new_n1927_) | ~new_n2040_ | ((new_n1931_ ^ ~P2_INSTADDRPOINTER_REG_13__SCAN_IN) & (new_n1797_ | new_n1927_)));
  assign new_n4432_ = (new_n2556_ | (P1_INSTADDRPOINTER_REG_16__SCAN_IN & ~new_n2522_ & new_n2552_) | (~P1_INSTADDRPOINTER_REG_16__SCAN_IN & (new_n2522_ | ~new_n2552_))) & new_n2596_ & (~new_n2556_ | (P1_INSTADDRPOINTER_REG_16__SCAN_IN ^ (~new_n2522_ & new_n2552_)));
  assign new_n4433_ = ~new_n4434_ & new_n4443_ & (new_n4441_ | ~new_n4449_) & (~new_n2596_ | (~new_n4436_ & ~new_n4438_ & new_n4439_));
  assign new_n4434_ = new_n4435_ & (((new_n2327_ | (~new_n2045_ & ~new_n2338_)) & (new_n2324_ | ~new_n2339_) & (~new_n2324_ | new_n2339_)) | ~new_n2503_ | (~new_n2327_ & (new_n2045_ | new_n2338_) & (new_n2324_ ^ new_n2339_)));
  assign new_n4435_ = (new_n2476_ | ~P1_EBX_REG_17__SCAN_IN) & (~new_n4027_ | ~new_n2476_ | ~new_n2053_);
  assign new_n4436_ = new_n4437_ & (~new_n2556_ | ~P1_INSTADDRPOINTER_REG_16__SCAN_IN) & ((~new_n2556_ & ~P1_INSTADDRPOINTER_REG_16__SCAN_IN) | (~new_n2522_ & new_n2552_));
  assign new_n4437_ = new_n2558_ ^ P1_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign new_n4438_ = ~new_n4437_ & ((new_n2556_ & P1_INSTADDRPOINTER_REG_16__SCAN_IN) | ((new_n2556_ | P1_INSTADDRPOINTER_REG_16__SCAN_IN) & (new_n2522_ | ~new_n2552_)));
  assign new_n4439_ = ~new_n4440_ ^ ((P1_INSTADDRPOINTER_REG_13__SCAN_IN & new_n2479_ & (new_n2310_ | ~new_n2047_ | new_n2244_) & (~new_n2310_ | (new_n2047_ & ~new_n2244_))) | ((P1_INSTADDRPOINTER_REG_13__SCAN_IN | (new_n2479_ & (new_n2310_ | ~new_n2047_ | new_n2244_) & (~new_n2310_ | (new_n2047_ & ~new_n2244_)))) & ((~new_n2680_ & (P1_INSTADDRPOINTER_REG_12__SCAN_IN | (new_n2479_ & (~new_n2047_ | new_n2244_) & (new_n2047_ | ~new_n2244_)))) | (P1_INSTADDRPOINTER_REG_12__SCAN_IN & new_n2479_ & (~new_n2047_ | new_n2244_) & (new_n2047_ | ~new_n2244_)))));
  assign new_n4440_ = ~P1_INSTADDRPOINTER_REG_14__SCAN_IN ^ (~new_n2479_ | (new_n2309_ & (new_n2311_ ^ new_n2163_)) | (~new_n2309_ & (new_n2311_ | ~new_n2163_) & (~new_n2311_ | new_n2163_)));
  assign new_n4441_ = (~new_n4442_ | (~new_n1648_ & ~new_n1696_) | ((~new_n1687_ | (new_n1649_ & ~new_n1697_)) & ~new_n1690_ & (~new_n1648_ | ~new_n1696_))) & new_n1758_ & (new_n4442_ | ((new_n1648_ | new_n1696_) & ((new_n1687_ & (~new_n1649_ | new_n1697_)) | new_n1690_ | (new_n1648_ & new_n1696_))));
  assign new_n4442_ = ~new_n1695_ & ~new_n1692_;
  assign new_n4443_ = ~new_n4444_ & (~new_n4448_ | ((~new_n4447_ | new_n2700_ | (new_n2695_ & ~new_n2701_)) & new_n2504_ & (new_n4447_ | (~new_n2700_ & (~new_n2695_ | new_n2701_)))));
  assign new_n4444_ = new_n4445_ & (~new_n2678_ | (new_n2671_ & (new_n1752_ | new_n1746_ | ~new_n1744_ | new_n1745_)) | (~new_n2671_ & ~new_n1752_ & ~new_n1746_ & new_n1744_ & ~new_n1745_));
  assign new_n4445_ = (new_n1759_ | ~P2_EAX_REG_31__SCAN_IN) & (~new_n4446_ | (new_n2976_ ? ~BUF1_REG_31__SCAN_IN : ~BUF2_REG_31__SCAN_IN));
  assign new_n4446_ = ~new_n1317_ & new_n1759_ & ~new_n1335_;
  assign new_n4447_ = ~new_n2321_ ^ (new_n2237_ & (~new_n2325_ | new_n2554_) & (new_n2325_ | ~new_n2554_));
  assign new_n4448_ = (new_n2505_ | ~P1_EAX_REG_15__SCAN_IN) & (~new_n2505_ | new_n2512_ | (~new_n2954_ & ~DATAI_15_) | (new_n2954_ & ~BUF1_REG_15__SCAN_IN));
  assign new_n4449_ = (~new_n1693_ | ~new_n2678_) & new_n4450_ & (~new_n4446_ | (new_n2976_ ? ~BUF1_REG_17__SCAN_IN : ~BUF2_REG_17__SCAN_IN));
  assign new_n4450_ = (new_n1759_ | ~P2_EAX_REG_17__SCAN_IN) & (~new_n1759_ | ~new_n1330_ | new_n1335_ | (new_n2976_ ? ~BUF1_REG_1__SCAN_IN : ~BUF2_REG_1__SCAN_IN));
  assign new_n4451_ = (new_n2045_ | new_n2327_ | new_n2338_) & new_n2504_ & (~new_n2045_ | (~new_n2327_ & ~new_n2338_));
  assign new_n4452_ = ((~new_n1637_ & new_n4454_) | ~new_n1758_ | (new_n1637_ & ~new_n4454_)) & new_n4458_ & ~new_n4456_ & ((new_n4455_ & (new_n4453_ | new_n4466_)) | ~new_n1758_ | (~new_n4455_ & ~new_n4453_ & ~new_n4466_));
  assign new_n4453_ = (new_n1641_ | (~new_n1647_ & new_n1698_)) & (new_n1700_ | (~new_n1699_ ^ ~new_n1486_));
  assign new_n4454_ = ~new_n1708_ & ~new_n1710_;
  assign new_n4455_ = ~new_n1638_ & ~new_n1640_;
  assign new_n4456_ = (new_n4457_ | (new_n2324_ & new_n2360_) | (~new_n2324_ & ~new_n2360_)) & (new_n2503_ | new_n2649_) & (~new_n4457_ | (new_n2324_ ^ new_n2360_));
  assign new_n4457_ = (~new_n2324_ | ~new_n2346_) & ((~new_n2324_ & ~new_n2346_) | ((~new_n2324_ | new_n2339_) & ((~new_n2324_ & new_n2339_) | (~new_n2327_ & (new_n2045_ | new_n2338_)))));
  assign new_n4458_ = ((new_n4459_ & ~P1_INSTADDRPOINTER_REG_21__SCAN_IN) | ~new_n2604_ | (~new_n4459_ & P1_INSTADDRPOINTER_REG_21__SCAN_IN)) & ((new_n4463_ & (~new_n2558_ ^ P1_INSTADDRPOINTER_REG_20__SCAN_IN)) | ~new_n2596_ | (~new_n4463_ & (~new_n2558_ | ~P1_INSTADDRPOINTER_REG_20__SCAN_IN) & (new_n2558_ | P1_INSTADDRPOINTER_REG_20__SCAN_IN)));
  assign new_n4459_ = (~new_n4461_ | new_n4460_ | (new_n2559_ & (~new_n2557_ | (~new_n2555_ & (new_n2522_ | ~new_n2552_))))) & (~new_n4462_ | ~new_n2559_ | (new_n2557_ & (new_n2555_ | (~new_n2522_ & new_n2552_))));
  assign new_n4460_ = new_n2558_ & P1_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign new_n4461_ = new_n2558_ & ~P1_INSTADDRPOINTER_REG_20__SCAN_IN & ~P1_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign new_n4462_ = ~new_n2558_ & (new_n2558_ | P1_INSTADDRPOINTER_REG_19__SCAN_IN) & (new_n2558_ | P1_INSTADDRPOINTER_REG_20__SCAN_IN);
  assign new_n4463_ = ~new_n4465_ & (new_n4464_ | (~new_n4460_ & (~new_n2559_ | (new_n2557_ & (new_n2555_ | (~new_n2522_ & new_n2552_))))));
  assign new_n4464_ = ~new_n2558_ & ~P1_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign new_n4465_ = new_n2558_ & P1_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign new_n4466_ = new_n1700_ & (~new_n1699_ | ~new_n1486_) & (new_n1699_ | new_n1486_);
  assign new_n4467_ = ((new_n2558_ & P1_INSTADDRPOINTER_REG_29__SCAN_IN) | (~new_n2558_ & ~P1_INSTADDRPOINTER_REG_29__SCAN_IN) | ((~new_n2558_ | new_n2612_) & (~new_n2558_ | new_n2617_) & ((~new_n2558_ & ~new_n2615_) | ~new_n2521_ | ~new_n2560_))) & new_n2604_ & ((new_n2558_ ^ P1_INSTADDRPOINTER_REG_29__SCAN_IN) | (new_n2558_ & ~new_n2612_) | (new_n2558_ & ~new_n2617_) | ((new_n2558_ | new_n2615_) & new_n2521_ & new_n2560_));
  assign new_n4468_ = ~new_n4469_ & (~new_n4473_ | (new_n2602_ & (~new_n2501_ | new_n2502_) & (new_n2501_ | ~new_n2502_))) & (~new_n2649_ | ((~new_n2501_ ^ ~new_n2502_) & (new_n2515_ ^ new_n2516_)));
  assign new_n4469_ = new_n4470_ & ((new_n4472_ & (~new_n1955_ | (new_n1952_ & (~new_n1951_ | (~new_n1796_ & new_n1937_))))) | ~new_n2040_ | (~new_n4472_ & new_n1955_ & (~new_n1952_ | (new_n1951_ & (new_n1796_ | ~new_n1937_)))));
  assign new_n4470_ = ((P2_INSTADDRPOINTER_REG_23__SCAN_IN & new_n1970_ & new_n1959_ & new_n1973_) | ~new_n2028_ | (~P2_INSTADDRPOINTER_REG_23__SCAN_IN & (~new_n1970_ | ~new_n1959_ | ~new_n1973_))) & new_n4471_ & (~new_n2682_ | ~new_n2004_);
  assign new_n4471_ = (~new_n2005_ | ~P2_PHYADDRPOINTER_REG_23__SCAN_IN) & (~P2_REIP_REG_23__SCAN_IN | new_n2005_ | ~new_n2022_) & (new_n2005_ | new_n2021_ | (new_n2730_ & P2_PHYADDRPOINTER_REG_23__SCAN_IN) | (~new_n2730_ & ~P2_PHYADDRPOINTER_REG_23__SCAN_IN));
  assign new_n4472_ = ~P2_INSTADDRPOINTER_REG_23__SCAN_IN ^ ((~new_n1947_ & (new_n1907_ | (new_n1330_ & P2_EBX_REG_23__SCAN_IN))) | new_n1534_ | (new_n1947_ & (~new_n1330_ | ~P2_EBX_REG_23__SCAN_IN)));
  assign new_n4473_ = new_n4474_ & (~new_n2604_ | (~new_n2656_ ^ (~new_n2561_ & (~new_n2521_ | ~new_n2560_))));
  assign new_n4474_ = (~new_n3502_ | ~P1_REIP_REG_23__SCAN_IN) & (~new_n2603_ | ~P1_PHYADDRPOINTER_REG_23__SCAN_IN) & (new_n2603_ | new_n3360_ | (~new_n2381_ & ~P1_PHYADDRPOINTER_REG_23__SCAN_IN) | (new_n2381_ & P1_PHYADDRPOINTER_REG_23__SCAN_IN));
  assign new_n4475_ = ~new_n4486_ & ~new_n4488_ & ~new_n4490_ & (~new_n4476_ | ((~new_n2039_ | (~new_n1795_ & P2_INSTADDRPOINTER_REG_25__SCAN_IN) | (new_n1795_ & ~P2_INSTADDRPOINTER_REG_25__SCAN_IN)) & new_n4420_ & (new_n2039_ | (~new_n1795_ ^ P2_INSTADDRPOINTER_REG_25__SCAN_IN))));
  assign new_n4476_ = new_n4477_ & (~new_n1526_ | ~new_n4485_) & ((P2_INSTADDRPOINTER_REG_25__SCAN_IN & new_n1958_ & P2_INSTADDRPOINTER_REG_23__SCAN_IN & P2_INSTADDRPOINTER_REG_24__SCAN_IN) | ~new_n2704_ | (~P2_INSTADDRPOINTER_REG_25__SCAN_IN & (~new_n1958_ | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN)));
  assign new_n4477_ = new_n4478_ & (~new_n4078_ | (new_n2003_ & (new_n2002_ | new_n2001_ | ~new_n1976_ | new_n2000_)) | (~new_n2003_ & ~new_n2002_ & ~new_n2001_ & new_n1976_ & ~new_n2000_));
  assign new_n4478_ = (~P2_REIP_REG_25__SCAN_IN | new_n4479_ | P2_STATE2_REG_2__SCAN_IN) & (~new_n4480_ | (new_n4482_ & P2_INSTADDRPOINTER_REG_25__SCAN_IN) | (~new_n4482_ & ~P2_INSTADDRPOINTER_REG_25__SCAN_IN)) & (~new_n4481_ | (new_n4484_ & P2_INSTADDRPOINTER_REG_25__SCAN_IN) | (~new_n4484_ & ~P2_INSTADDRPOINTER_REG_25__SCAN_IN)) & (~new_n4479_ | ~P2_INSTADDRPOINTER_REG_25__SCAN_IN);
  assign new_n4479_ = ~new_n2706_ & ~new_n4031_;
  assign new_n4480_ = new_n2706_ & new_n1783_;
  assign new_n4481_ = new_n2706_ & ~new_n4055_;
  assign new_n4482_ = new_n4483_ & new_n4063_;
  assign new_n4483_ = new_n1971_ & new_n1969_ & new_n1973_ & new_n1972_ & P2_INSTADDRPOINTER_REG_7__SCAN_IN & P2_INSTADDRPOINTER_REG_8__SCAN_IN & P2_INSTADDRPOINTER_REG_23__SCAN_IN & P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign new_n4484_ = new_n4483_ & P2_INSTADDRPOINTER_REG_6__SCAN_IN & P2_INSTADDRPOINTER_REG_5__SCAN_IN & P2_INSTADDRPOINTER_REG_3__SCAN_IN & P2_INSTADDRPOINTER_REG_4__SCAN_IN & P2_INSTADDRPOINTER_REG_2__SCAN_IN & P2_INSTADDRPOINTER_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign new_n4485_ = new_n2706_ & (new_n2667_ | new_n2684_ | (new_n1787_ & new_n1764_));
  assign new_n4486_ = new_n4487_ & (((~new_n2368_ | (~new_n2501_ & new_n2423_)) & (~new_n2324_ | new_n2419_) & (new_n2324_ | ~new_n2419_)) | ~new_n2503_ | (new_n2368_ & (new_n2501_ | ~new_n2423_) & (~new_n2324_ ^ ~new_n2419_)));
  assign new_n4487_ = (new_n2476_ | ~P1_EBX_REG_25__SCAN_IN) & ((~new_n2451_ & (new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_25__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_25__SCAN_IN)))) | ~new_n2476_ | ~new_n2053_ | (new_n2451_ & (new_n2090_ | (new_n2456_ & P1_INSTADDRPOINTER_REG_25__SCAN_IN) | (~new_n2455_ & P1_EBX_REG_25__SCAN_IN)) & (~new_n2090_ | ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_25__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_25__SCAN_IN)))));
  assign new_n4488_ = new_n4489_ & (((new_n2324_ ^ new_n2382_) & (~new_n2324_ | ~new_n2369_) & (new_n2501_ | (~new_n2324_ & ~new_n2369_))) | ~new_n2504_ | ((new_n2324_ | ~new_n2382_) & (~new_n2324_ | new_n2382_) & ((new_n2324_ & new_n2369_) | (~new_n2501_ & (new_n2324_ | new_n2369_)))));
  assign new_n4489_ = (~new_n2505_ | ~new_n2513_ | (new_n2954_ & ~BUF1_REG_8__SCAN_IN) | (~new_n2954_ & ~DATAI_8_)) & (new_n3230_ | ~new_n2505_ | ~new_n2291_) & (new_n2505_ | ~P1_EAX_REG_24__SCAN_IN);
  assign new_n4490_ = new_n2602_ & (new_n2439_ ^ (~new_n2043_ & ~new_n2449_));
  assign new_n4491_ = ~new_n4493_ & (~new_n4504_ | ((~new_n4492_ | (~new_n1306_ & (~new_n1526_ | (new_n1308_ & new_n1630_) | (~new_n1308_ & ~new_n1630_)))) & new_n1758_ & (new_n4492_ | new_n1306_ | (new_n1526_ & (~new_n1308_ | ~new_n1630_) & (new_n1308_ | new_n1630_)))));
  assign new_n4492_ = ~new_n1728_ & ~new_n1712_;
  assign new_n4493_ = new_n4502_ & ((((new_n2324_ | new_n2440_) & ~new_n2043_ & ~new_n2449_) ? (~new_n4503_ & (new_n2324_ | ~new_n4494_)) : ((~new_n2324_ | new_n4494_) & new_n4503_ & (~new_n2324_ | ~new_n2440_))) | ~new_n4501_ | (~new_n4503_ & new_n2324_ & ~new_n4494_) | (~new_n4503_ & new_n2324_ & new_n2440_) | (new_n4503_ & ~new_n2324_ & new_n4494_));
  assign new_n4494_ = (new_n4495_ | (~P1_STATEBS16_REG_SCAN_IN & ~P1_STATE2_REG_2__SCAN_IN)) & ((~P1_PHYADDRPOINTER_REG_30__SCAN_IN & (P1_STATEBS16_REG_SCAN_IN | (P1_PHYADDRPOINTER_REG_29__SCAN_IN & P1_PHYADDRPOINTER_REG_28__SCAN_IN & new_n2418_ & P1_PHYADDRPOINTER_REG_27__SCAN_IN))) | P1_STATE2_REG_2__SCAN_IN | (P1_PHYADDRPOINTER_REG_30__SCAN_IN & ~P1_STATEBS16_REG_SCAN_IN & (~P1_PHYADDRPOINTER_REG_29__SCAN_IN | ~P1_PHYADDRPOINTER_REG_28__SCAN_IN | ~new_n2418_ | ~P1_PHYADDRPOINTER_REG_27__SCAN_IN)));
  assign new_n4495_ = (~new_n2292_ | ~P1_EAX_REG_30__SCAN_IN) & ((~new_n4496_ & (~new_n2331_ | (new_n2442_ & new_n2443_))) | ~new_n2237_ | (new_n4496_ & (~new_n2442_ | ~new_n2443_)));
  assign new_n4496_ = new_n4497_ & new_n4498_ & new_n4500_ & (~new_n2056_ | ~P1_INSTQUEUE_REG_3__7__SCAN_IN) & (~new_n2099_ | ~P1_INSTQUEUE_REG_7__7__SCAN_IN);
  assign new_n4497_ = (~new_n2098_ | ~P1_INSTQUEUE_REG_10__7__SCAN_IN) & (~new_n2057_ | ~P1_INSTQUEUE_REG_15__7__SCAN_IN) & (~new_n2080_ | ~P1_INSTQUEUE_REG_11__7__SCAN_IN);
  assign new_n4498_ = new_n4499_ & (~P1_INSTQUEUE_REG_0__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_1__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_14__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  assign new_n4499_ = (~P1_INSTQUEUE_REG_2__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_13__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_12__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_4__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n4500_ = (~P1_INSTQUEUE_REG_9__7__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_6__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN) & (~P1_INSTQUEUE_REG_8__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN) & (~P1_INSTQUEUE_REG_5__7__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  assign new_n4501_ = new_n2505_ & new_n2053_;
  assign new_n4502_ = (new_n2505_ | ~P1_EAX_REG_31__SCAN_IN) & (~new_n2505_ | ~new_n2291_ | (new_n2954_ ? ~BUF1_REG_31__SCAN_IN : ~DATAI_31_));
  assign new_n4503_ = (~P1_PHYADDRPOINTER_REG_31__SCAN_IN | ~P1_STATEBS16_REG_SCAN_IN | P1_STATE2_REG_2__SCAN_IN) & (~P1_EAX_REG_31__SCAN_IN | ~new_n2053_ | ~P1_STATE2_REG_2__SCAN_IN) & (~new_n2644_ | P1_STATEBS16_REG_SCAN_IN | P1_STATE2_REG_2__SCAN_IN);
  assign new_n4504_ = (~new_n1713_ | ~new_n2678_) & new_n4505_ & (~new_n4446_ | (new_n2976_ ? ~BUF1_REG_26__SCAN_IN : ~BUF2_REG_26__SCAN_IN));
  assign new_n4505_ = (new_n1759_ | ~P2_EAX_REG_26__SCAN_IN) & (~new_n1759_ | ~new_n1330_ | new_n1335_ | (new_n2976_ ? ~BUF1_REG_10__SCAN_IN : ~BUF2_REG_10__SCAN_IN));
  assign new_n4506_ = new_n4507_ & (((~new_n2324_ | new_n2414_) & (new_n2324_ | ~new_n2414_) & (new_n2324_ | ~new_n2419_) & ((~new_n2501_ & new_n2423_) | ~new_n2368_ | (new_n2324_ & ~new_n2419_))) | ~new_n2503_ | ((~new_n2324_ ^ ~new_n2414_) & ((~new_n2324_ & new_n2419_) | ((new_n2501_ | ~new_n2423_) & new_n2368_ & (~new_n2324_ | new_n2419_)))));
  assign new_n4507_ = (new_n2476_ | ~P1_EBX_REG_26__SCAN_IN) & ((~new_n2450_ & (~new_n2090_ | (new_n2456_ & P1_INSTADDRPOINTER_REG_26__SCAN_IN) | (~new_n2455_ & P1_EBX_REG_26__SCAN_IN)) & (new_n2090_ | ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_26__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_26__SCAN_IN)))) | ~new_n2476_ | ~new_n2053_ | (new_n2450_ & (~new_n2090_ ^ ((~new_n2456_ | ~P1_INSTADDRPOINTER_REG_26__SCAN_IN) & (new_n2455_ | ~P1_EBX_REG_26__SCAN_IN)))));
  assign new_n4508_ = (new_n2031_ | P2_INSTADDRPOINTER_REG_29__SCAN_IN) & ((new_n2031_ & P2_INSTADDRPOINTER_REG_29__SCAN_IN) | ~new_n2038_ | ((new_n2039_ | (~new_n1795_ & P2_INSTADDRPOINTER_REG_25__SCAN_IN)) & new_n2034_ & (~new_n1795_ | P2_INSTADDRPOINTER_REG_25__SCAN_IN)));
  assign new_n4509_ = new_n4510_ & ((P2_INSTADDRPOINTER_REG_30__SCAN_IN & new_n2029_ & P2_INSTADDRPOINTER_REG_29__SCAN_IN & new_n1958_ & P2_INSTADDRPOINTER_REG_23__SCAN_IN & P2_INSTADDRPOINTER_REG_24__SCAN_IN) | ~new_n2704_ | (~P2_INSTADDRPOINTER_REG_30__SCAN_IN & (~new_n2029_ | ~P2_INSTADDRPOINTER_REG_29__SCAN_IN | ~new_n1958_ | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN)));
  assign new_n4510_ = (~new_n1751_ | ~new_n4485_) & new_n4511_ & ((new_n2689_ & ~new_n2692_) | ~new_n4078_ | (~new_n2689_ & new_n2692_));
  assign new_n4511_ = new_n4512_ & (~P2_REIP_REG_30__SCAN_IN | new_n4479_ | P2_STATE2_REG_2__SCAN_IN);
  assign new_n4512_ = (~new_n4480_ | (P2_INSTADDRPOINTER_REG_30__SCAN_IN & new_n4482_ & new_n4513_) | (~P2_INSTADDRPOINTER_REG_30__SCAN_IN & (~new_n4482_ | ~new_n4513_))) & (~new_n4479_ | ~P2_INSTADDRPOINTER_REG_30__SCAN_IN) & (~new_n4481_ | (~P2_INSTADDRPOINTER_REG_30__SCAN_IN ^ (new_n4484_ & new_n4513_)));
  assign new_n4513_ = new_n2029_ & P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign new_n4514_ = (new_n2773_ | (~new_n1907_ & (~new_n1330_ | ~P2_EBX_REG_30__SCAN_IN))) & ~new_n1534_ & (~new_n2773_ | new_n1907_ | (new_n1330_ & P2_EBX_REG_30__SCAN_IN));
endmodule


