// Benchmark "multiplier_15_sat" written by ABC on Mon Nov 14 17:45:49 2022

module multiplier_15_sat ( 
    \a[0] , \a[1] , \a[2] , \b[0] , \b[1] ,
    sat  );
  input  \a[0] , \a[1] , \a[2] , \b[0] , \b[1] ;
  output sat;
  assign sat = ((~\a[2]  | \b[1] ) ^ ((\a[2]  & \b[0]  & ((\a[0]  ? ~\b[0]  : \a[1] ) | ~\b[1]  | (~\a[1]  ^ \a[2] ))) | ((((\a[0]  ? \b[0]  : ~\a[1] ) & \b[1]  & (\a[1]  ^ \a[2] )) ^ (\a[2]  & ~\b[0] )) & (~\b[1]  | ((\a[0]  | ~\a[1] ) & ((~\a[1]  ^ \a[2] ) | ~\a[0]  | (\b[0]  & \b[1] )))) & ((~\a[1]  ^ \a[2] ) | ~\a[0]  | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & (~\b[0]  | \a[0]  | ~\a[1] ) & ((~\a[1]  & \a[2] ) | (\a[1]  & ~\a[2] ) | ~\a[0]  | ~\b[1] ) & (~\a[2]  | ~\b[0]  | \a[0]  | \a[1] ) & \a[2]  & (~\a[0]  | ~\b[0] )))) & ((~\a[1]  ^ \a[2] ) | ~\a[0]  | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & (~\b[0]  | \a[0]  | ~\a[1] ) & ((~\a[1]  & \a[2] ) | (\a[1]  & ~\a[2] ) | ~\a[0]  | ~\b[1] ) & ~\a[1]  & \a[2]  & \b[0]  & \a[0]  & \b[1] ;
endmodule


