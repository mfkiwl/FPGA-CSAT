// Benchmark "multiplier_9991_sat" written by ABC on Fri Nov 11 15:23:58 2022

module multiplier_9991_sat ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] ,
    sat  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \b[0] , \b[1] , \b[2] ,
    \b[3] , \b[4] , \b[5] , \b[6] ;
  output sat;
  wire new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_,
    new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_,
    new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_,
    new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_,
    new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_;
  assign sat = (new_n24_ | (\a[2]  & (new_n25_ | ~new_n100_) & (~new_n25_ | new_n100_)) | (((new_n101_ & \a[2] ) | ((~new_n101_ | ~\a[2] ) & (new_n101_ | \a[2] ) & ((new_n102_ & \a[2] ) | (~new_n103_ & (~new_n102_ | ~\a[2] ) & (new_n102_ | \a[2] ))))) & (~\a[2]  | (~new_n25_ & new_n100_) | (new_n25_ & ~new_n100_)) & (\a[2]  | (~new_n25_ ^ new_n100_)))) & new_n99_ & (~new_n24_ | ((~\a[2]  | (~new_n25_ & new_n100_) | (new_n25_ & ~new_n100_)) & (((~new_n101_ | ~\a[2] ) & ((new_n101_ & \a[2] ) | (~new_n101_ & ~\a[2] ) | ((~new_n102_ | ~\a[2] ) & (new_n103_ | (new_n102_ & \a[2] ) | (~new_n102_ & ~\a[2] ))))) | (\a[2]  & (new_n25_ | ~new_n100_) & (~new_n25_ | new_n100_)) | (~\a[2]  & (new_n25_ ^ new_n100_)))));
  assign new_n24_ = new_n98_ ^ (((\a[5]  & (((~new_n65_ | ~\a[8] ) & (new_n95_ | (new_n65_ & \a[8] ) | (~new_n65_ & ~\a[8] ))) | (new_n96_ & \a[8] ) | (~new_n96_ & ~\a[8] )) & ((new_n65_ & \a[8] ) | (~new_n95_ & (~new_n65_ | ~\a[8] ) & (new_n65_ | \a[8] )) | (new_n96_ ^ \a[8] ))) | (~new_n25_ & (~\a[5]  | (((new_n65_ & \a[8] ) | (~new_n95_ & (~new_n65_ | ~\a[8] ) & (new_n65_ | \a[8] ))) & (~new_n96_ | ~\a[8] ) & (new_n96_ | \a[8] )) | ((~new_n65_ | ~\a[8] ) & (new_n95_ | (new_n65_ & \a[8] ) | (~new_n65_ & ~\a[8] )) & (~new_n96_ ^ \a[8] ))) & (\a[5]  | (((new_n65_ & \a[8] ) | (~new_n95_ & (~new_n65_ | ~\a[8] ) & (new_n65_ | \a[8] ))) ^ (new_n96_ ^ \a[8] ))))) ^ (~new_n92_ ^ (\a[8]  ^ ((new_n96_ & \a[8] ) | (((new_n65_ & \a[8] ) | (~new_n95_ & (~new_n65_ | ~\a[8] ) & (new_n65_ | \a[8] ))) & (~new_n96_ | ~\a[8] ) & (new_n96_ | \a[8] ))))));
  assign new_n25_ = (~new_n26_ | ~\a[5] ) & ((new_n26_ & \a[5] ) | (~new_n26_ & ~\a[5] ) | ((~new_n71_ | ~\a[5] ) & ((new_n71_ & \a[5] ) | (~new_n71_ & ~\a[5] ) | ((~new_n72_ | ~\a[5] ) & (((~\a[5]  | (~new_n48_ & new_n64_) | (new_n48_ & ~new_n64_)) & (new_n73_ | (\a[5]  & (new_n48_ | ~new_n64_) & (~new_n48_ | new_n64_)) | (~\a[5]  & (new_n48_ ^ new_n64_)))) | (new_n72_ & \a[5] ) | (~new_n72_ & ~\a[5] ))))));
  assign new_n26_ = (new_n65_ ^ \a[8] ) ^ ((\a[8]  & (new_n27_ | ~new_n68_) & (~new_n27_ | new_n68_)) | (((new_n44_ & \a[8] ) | ((new_n45_ | (~new_n48_ & new_n64_)) & (~new_n44_ | ~\a[8] ) & (new_n44_ | \a[8] ))) & (~\a[8]  | (~new_n27_ & new_n68_) | (new_n27_ & ~new_n68_)) & (\a[8]  | (~new_n27_ ^ new_n68_))));
  assign new_n27_ = ~new_n28_ & (~new_n43_ | (~new_n32_ & (new_n35_ | ~new_n42_)));
  assign new_n28_ = (~\a[11]  ^ (new_n31_ & (~new_n29_ | ~new_n30_))) & ((\b[3]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] )) | (\b[2]  & \a[11]  & \a[12] ));
  assign new_n29_ = (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] );
  assign new_n30_ = ((\b[4]  & \b[5] ) | (((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))) & (~\b[4]  | ~\b[5] ) & (\b[4]  | \b[5] ))) ^ (\b[5]  ^ \b[6] );
  assign new_n31_ = (~\b[4]  | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\a[8]  ^ \a[9] ) | (~\a[9]  ^ ~\a[10] )) & (~\b[5]  | (\a[8]  ^ \a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[6]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  ^ ~\a[11] ));
  assign new_n32_ = (~\a[11]  ^ (new_n34_ & (~new_n29_ | ~new_n33_))) & ((\b[2]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] )) | (\b[1]  & \a[11]  & \a[12] ));
  assign new_n33_ = ((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))) ^ (\b[4]  ^ \b[5] );
  assign new_n34_ = (~\b[3]  | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\a[8]  ^ \a[9] ) | (~\a[9]  ^ ~\a[10] )) & (~\b[4]  | (\a[8]  ^ \a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[5]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  ^ ~\a[11] ));
  assign new_n35_ = (new_n38_ | (\a[11]  ^ (new_n37_ & (~new_n29_ | ~new_n36_)))) & ((~new_n39_ & (new_n40_ | ~new_n41_)) | (~new_n38_ & (~\a[11]  ^ (new_n37_ & (~new_n29_ | ~new_n36_)))) | (new_n38_ & (~\a[11]  | ~new_n37_ | (new_n29_ & new_n36_)) & (\a[11]  | (new_n37_ & (~new_n29_ | ~new_n36_)))));
  assign new_n36_ = (\b[3]  ^ \b[4] ) ^ ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] )));
  assign new_n37_ = (~\b[2]  | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\a[8]  ^ \a[9] ) | (~\a[9]  ^ ~\a[10] )) & (~\b[3]  | (\a[8]  ^ \a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[4]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  ^ ~\a[11] ));
  assign new_n38_ = (~\b[1]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] )) & (~\b[0]  | ~\a[11]  | ~\a[12] );
  assign new_n39_ = \b[0]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] ) & (~\b[0]  | (\a[8]  ^ \a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[11]  & (~\b[0]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] )) & (~\b[0]  | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\a[8]  ^ \a[9] ) | (~\a[9]  ^ ~\a[10] )) & ((\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[1]  | (\a[8]  ^ \a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ));
  assign new_n40_ = \a[11]  ^ (((\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\a[8]  ^ \a[9] ) | (~\a[9]  ^ ~\a[10] )) & (~\b[3]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[2]  | (\a[8]  ^ \a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )));
  assign new_n41_ = (\b[0]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] )) ^ ((~\b[0]  | (\a[8]  ^ \a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[11]  & (~\b[0]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] )) & (~\b[0]  | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\a[8]  ^ \a[9] ) | (~\a[9]  ^ ~\a[10] )) & ((\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  ^ ~\a[11] )) & (~\b[1]  | (\a[8]  ^ \a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )));
  assign new_n42_ = (~\a[11]  ^ (new_n34_ & (~new_n29_ | ~new_n33_))) ^ ((\b[2]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] )) | (\b[1]  & \a[11]  & \a[12] ));
  assign new_n43_ = (~\a[11]  ^ (new_n31_ & (~new_n29_ | ~new_n30_))) ^ ((\b[3]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] )) | (\b[2]  & \a[11]  & \a[12] ));
  assign new_n44_ = new_n43_ ^ (new_n32_ | (~new_n35_ & new_n42_));
  assign new_n45_ = ~new_n46_ & (new_n35_ | ~new_n42_) & (~new_n35_ | new_n42_);
  assign new_n46_ = \a[8]  ^ (~\b[6]  | ((new_n47_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] ))));
  assign new_n47_ = (~\b[5]  | ~\b[6] ) & (((~\b[4]  | ~\b[5] ) & (((~\b[3]  | ~\b[4] ) & ((\b[3]  & \b[4] ) | (~\b[3]  & ~\b[4] ) | ((~\b[2]  | ~\b[3] ) & ((~\b[2]  & ~\b[3] ) | (\b[2]  & \b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] ))))) | (\b[4]  & \b[5] ) | (~\b[4]  & ~\b[5] ))) | (\b[5]  & \b[6] ) | (~\b[5]  & ~\b[6] ));
  assign new_n48_ = (new_n51_ | (~new_n49_ & new_n50_) | (new_n49_ & ~new_n50_)) & (((~new_n52_ | new_n53_) & (((new_n54_ | ~new_n63_) & (new_n57_ | (~new_n54_ & new_n63_) | (new_n54_ & ~new_n63_))) | (~new_n52_ & new_n53_) | (new_n52_ & ~new_n53_))) | (~new_n51_ & (new_n49_ | ~new_n50_) & (~new_n49_ | new_n50_)) | (new_n51_ & (new_n49_ ^ new_n50_)));
  assign new_n49_ = ~new_n39_ & (new_n40_ | ~new_n41_);
  assign new_n50_ = ~new_n38_ ^ (~\a[11]  ^ (new_n37_ & (~new_n29_ | ~new_n36_)));
  assign new_n51_ = \a[8]  ^ (((new_n47_ ^ \b[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[5]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[6]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n52_ = ~new_n40_ ^ new_n41_;
  assign new_n53_ = \a[8]  ^ ((~new_n30_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[4]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[5]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[6]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )));
  assign new_n54_ = \a[8]  ^ (new_n56_ & (~new_n33_ | ~new_n55_));
  assign new_n55_ = (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] );
  assign new_n56_ = (~\b[4]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[5]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[3]  | (~\a[6]  ^ ~\a[7] ) | (\a[5]  ^ \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ));
  assign new_n57_ = (~new_n59_ | (\a[8]  ^ (new_n58_ & (~new_n36_ | ~new_n55_)))) & ((~new_n60_ & (new_n61_ | ~new_n62_)) | (new_n59_ & (~\a[8]  ^ (new_n58_ & (~new_n36_ | ~new_n55_)))) | (~new_n59_ & (~\a[8]  | ~new_n58_ | (new_n36_ & new_n55_)) & (\a[8]  | (new_n58_ & (~new_n36_ | ~new_n55_)))));
  assign new_n58_ = (~\b[3]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[4]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[2]  | (~\a[6]  ^ ~\a[7] ) | (\a[5]  ^ \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ));
  assign new_n59_ = ((\b[0]  & (~\a[8]  ^ \a[9] ) & (\a[9]  | \a[10] ) & (~\a[9]  | ~\a[10] )) | (\b[1]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] ) & (\a[10]  ^ ~\a[11] )) | ((~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[11]  & \b[0]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] ));
  assign new_n60_ = \b[0]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] ) & (~\b[0]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[8]  & (~\b[0]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] )) & ((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[1]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (\a[5]  ^ \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ));
  assign new_n61_ = \a[8]  ^ (((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[2]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[6]  ^ ~\a[7] ) | (\a[5]  ^ \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )));
  assign new_n62_ = (\b[0]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] )) ^ ((~\b[0]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[8]  & (~\b[0]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] )) & ((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[1]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (\a[5]  ^ \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )));
  assign new_n63_ = ((~\b[0]  | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\a[8]  ^ \a[9] ) | (~\a[9]  ^ ~\a[10] )) & (~\b[1]  | (\a[8]  ^ \a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[2]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))) ^ (~\a[11]  | ((~\b[0]  | (\a[8]  ^ \a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[11]  & (~\b[0]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ))));
  assign new_n64_ = ~new_n46_ ^ (~new_n35_ ^ new_n42_);
  assign new_n65_ = new_n69_ ^ (new_n66_ | (new_n68_ & (new_n28_ | (new_n43_ & (new_n32_ | (~new_n35_ & new_n42_))))));
  assign new_n66_ = ~new_n67_ & (~\a[11]  ^ (((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~new_n47_ ^ ~\b[6] )) & (~\b[5]  | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\a[9]  ^ \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[6]  | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] ) | (~\a[8]  ^ ~\a[9] ))));
  assign new_n67_ = (~\b[4]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] )) & (~\b[3]  | ~\a[11]  | ~\a[12] );
  assign new_n68_ = ~new_n67_ ^ (~\a[11]  ^ (((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~new_n47_ ^ ~\b[6] )) & (~\b[5]  | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\a[9]  ^ \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[6]  | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] ) | (~\a[8]  ^ ~\a[9] ))));
  assign new_n69_ = ((\b[5]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] )) | (\b[4]  & \a[11]  & \a[12] )) ^ (~\a[11]  ^ (~\b[6]  | (~new_n70_ & (~new_n29_ | new_n47_))));
  assign new_n70_ = (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] ) & (~\a[8]  ^ \a[9] ) & (\a[9]  ^ ~\a[10] );
  assign new_n71_ = ((new_n44_ & \a[8] ) | ((~new_n44_ | ~\a[8] ) & (new_n44_ | \a[8] ) & (new_n45_ | (~new_n48_ & new_n64_)))) ^ (\a[8]  ^ (~new_n27_ ^ new_n68_));
  assign new_n72_ = (new_n45_ | (~new_n48_ & new_n64_)) ^ (new_n44_ ^ \a[8] );
  assign new_n73_ = (~new_n75_ | ~\a[5] ) & ((new_n75_ & \a[5] ) | (~new_n75_ & ~\a[5] ) | ((~\a[5]  | (new_n74_ & ((~new_n54_ & new_n63_) | (~new_n57_ & (new_n54_ | ~new_n63_) & (~new_n54_ | new_n63_)))) | (~new_n74_ & (new_n54_ | ~new_n63_) & (new_n57_ | (~new_n54_ & new_n63_) | (new_n54_ & ~new_n63_)))) & ((\a[5]  & (~new_n74_ | ((new_n54_ | ~new_n63_) & (new_n57_ | (~new_n54_ & new_n63_) | (new_n54_ & ~new_n63_)))) & (new_n74_ | (~new_n54_ & new_n63_) | (~new_n57_ & (new_n54_ | ~new_n63_) & (~new_n54_ | new_n63_)))) | (~\a[5]  & (~new_n74_ ^ ((~new_n54_ & new_n63_) | (~new_n57_ & (new_n54_ | ~new_n63_) & (~new_n54_ | new_n63_))))) | ((new_n91_ | (~new_n57_ & (new_n54_ | ~new_n63_) & (~new_n54_ | new_n63_)) | (new_n57_ & (new_n54_ ^ new_n63_))) & (new_n76_ | (~new_n91_ & (new_n57_ | (~new_n54_ & new_n63_) | (new_n54_ & ~new_n63_)) & (~new_n57_ | (~new_n54_ ^ new_n63_))) | (new_n91_ & (new_n57_ ^ (~new_n54_ ^ new_n63_))))))));
  assign new_n74_ = ~new_n52_ ^ new_n53_;
  assign new_n75_ = ((new_n52_ & ~new_n53_) | (((~new_n54_ & new_n63_) | (~new_n57_ & (new_n54_ | ~new_n63_) & (~new_n54_ | new_n63_))) & (new_n52_ | ~new_n53_) & (~new_n52_ | new_n53_))) ^ (~new_n51_ ^ (~new_n49_ ^ new_n50_));
  assign new_n76_ = (~new_n77_ | new_n78_) & ((~new_n77_ & new_n78_) | (new_n77_ & ~new_n78_) | ((~new_n79_ | new_n80_) & ((~new_n79_ & new_n80_) | (new_n79_ & ~new_n80_) | ((new_n81_ | ~new_n90_) & (new_n84_ | (~new_n81_ & new_n90_) | (new_n81_ & ~new_n90_))))));
  assign new_n77_ = (new_n60_ | (~new_n61_ & new_n62_)) ^ (new_n59_ ^ (~\a[8]  ^ (new_n58_ & (~new_n36_ | ~new_n55_))));
  assign new_n78_ = \a[5]  ^ (((new_n47_ ^ \b[6] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[5]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[6]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n79_ = ~new_n61_ ^ new_n62_;
  assign new_n80_ = \a[5]  ^ ((~new_n30_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[4]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[5]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[6]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )));
  assign new_n81_ = \a[5]  ^ (new_n83_ & (~new_n33_ | ~new_n82_));
  assign new_n82_ = (~\a[2]  | ~\a[3] ) & (\a[2]  | \a[3] ) & (\a[4]  | \a[5] ) & (~\a[4]  | ~\a[5] );
  assign new_n83_ = (~\b[4]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[5]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[3]  | (~\a[3]  ^ ~\a[4] ) | (\a[2]  ^ \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n84_ = (~new_n86_ | (\a[5]  ^ (new_n85_ & (~new_n36_ | ~new_n82_)))) & ((~new_n87_ & (new_n88_ | ~new_n89_)) | (new_n86_ & (~\a[5]  ^ (new_n85_ & (~new_n36_ | ~new_n82_)))) | (~new_n86_ & (~\a[5]  | ~new_n85_ | (new_n36_ & new_n82_)) & (\a[5]  | (new_n85_ & (~new_n36_ | ~new_n82_)))));
  assign new_n85_ = (~\b[3]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[4]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[2]  | (~\a[3]  ^ ~\a[4] ) | (\a[2]  ^ \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n86_ = ((\b[0]  & (~\a[5]  ^ \a[6] ) & (\a[6]  | \a[7] ) & (~\a[6]  | ~\a[7] )) | (\b[1]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  ^ ~\a[8] )) | ((~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[8]  & \b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ));
  assign new_n87_ = \b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (~\b[0]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[5]  & (~\b[0]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] )) & ((\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[1]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (\a[2]  ^ \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n88_ = \a[5]  ^ (((\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[2]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[3]  ^ ~\a[4] ) | (\a[2]  ^ \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )));
  assign new_n89_ = (\b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] )) ^ ((~\b[0]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[5]  & (~\b[0]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] )) & ((\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[1]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (\a[2]  ^ \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )));
  assign new_n90_ = (~\a[8]  | ((~\b[0]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[8]  & (~\b[0]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] )))) ^ ((~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (\a[5]  ^ \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )) & (~\b[1]  | (\a[5]  ^ \a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[2]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n91_ = \a[5]  ^ (~\b[6]  | ((new_n47_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] ))));
  assign new_n92_ = (~\a[11]  | ((~\b[6]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] )) & (~\a[12]  | ~\b[5] ))) & ((~new_n94_ & (new_n93_ | ~new_n69_)) | (\a[11]  & ((\b[6]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] )) | (\a[12]  & \b[5] ))) | (~\a[11]  & (~\a[12]  | ~\b[6] )));
  assign new_n93_ = ~new_n66_ & (new_n27_ | ~new_n68_);
  assign new_n94_ = ((\b[5]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] )) | (\b[4]  & \a[11]  & \a[12] )) & (~\a[11]  ^ (~\b[6]  | (~new_n70_ & (~new_n29_ | new_n47_))));
  assign new_n95_ = (~\a[8]  | (~new_n27_ & new_n68_) | (new_n27_ & ~new_n68_)) & (((~new_n44_ | ~\a[8] ) & ((new_n44_ & \a[8] ) | (~new_n44_ & ~\a[8] ) | (~new_n45_ & (new_n48_ | ~new_n64_)))) | (\a[8]  & (new_n27_ | ~new_n68_) & (~new_n27_ | new_n68_)) | (~\a[8]  & (new_n27_ ^ new_n68_)));
  assign new_n96_ = new_n97_ ^ (new_n94_ | (new_n69_ & (new_n66_ | (~new_n27_ & new_n68_))));
  assign new_n97_ = \a[11]  ? ((~\a[12]  | ~\b[5] ) & (~\b[6]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ))) : (\a[12]  & \b[6] );
  assign new_n98_ = \a[2]  ^ (~\a[5]  ^ (\a[11]  & (~\a[12]  | ~\b[6] )));
  assign new_n99_ = ((~\a[2]  ^ (~new_n25_ ^ new_n100_)) ^ ((new_n101_ & \a[2] ) | ((~new_n101_ | ~\a[2] ) & (new_n101_ | \a[2] ) & ((new_n102_ & \a[2] ) | (~new_n103_ & (~new_n102_ | ~\a[2] ) & (new_n102_ | \a[2] )))))) & ((~new_n101_ ^ \a[2] ) ^ ((new_n102_ & \a[2] ) | (~new_n103_ & (~new_n102_ | ~\a[2] ) & (new_n102_ | \a[2] )))) & ~new_n128_ & new_n129_ & (new_n103_ ^ (new_n102_ ^ \a[2] ));
  assign new_n100_ = \a[5]  ^ (((new_n65_ & \a[8] ) | (~new_n95_ & (~new_n65_ | ~\a[8] ) & (new_n65_ | \a[8] ))) ^ (new_n96_ ^ \a[8] ));
  assign new_n101_ = (new_n26_ ^ \a[5] ) ^ ((new_n71_ & \a[5] ) | ((~new_n71_ | ~\a[5] ) & (new_n71_ | \a[5] ) & ((new_n72_ & \a[5] ) | (((\a[5]  & (new_n48_ | ~new_n64_) & (~new_n48_ | new_n64_)) | (~new_n73_ & (~\a[5]  | (~new_n48_ & new_n64_) | (new_n48_ & ~new_n64_)) & (\a[5]  | (~new_n48_ ^ new_n64_)))) & (~new_n72_ | ~\a[5] ) & (new_n72_ | \a[5] )))));
  assign new_n102_ = ((new_n72_ & \a[5] ) | (((\a[5]  & (new_n48_ | ~new_n64_) & (~new_n48_ | new_n64_)) | (~new_n73_ & (~\a[5]  | (~new_n48_ & new_n64_) | (new_n48_ & ~new_n64_)) & (\a[5]  | (~new_n48_ ^ new_n64_)))) & (~new_n72_ | ~\a[5] ) & (new_n72_ | \a[5] ))) ^ (new_n71_ ^ \a[5] );
  assign new_n103_ = (~\a[2]  | ((~new_n72_ | ~\a[5] ) & (new_n72_ | \a[5] ) & ((new_n104_ & \a[5] ) | (~new_n73_ & (~new_n104_ | ~\a[5] ) & (new_n104_ | \a[5] )))) | ((~new_n72_ ^ \a[5] ) & (~new_n104_ | ~\a[5] ) & (new_n73_ | (new_n104_ & \a[5] ) | (~new_n104_ & ~\a[5] )))) & (((~\a[2]  | (~new_n73_ & (~new_n104_ | ~\a[5] ) & (new_n104_ | \a[5] )) | (new_n73_ & (~new_n104_ ^ \a[5] ))) & (((~new_n105_ | ~\a[2] ) & (new_n106_ | (new_n105_ & \a[2] ) | (~new_n105_ & ~\a[2] ))) | (\a[2]  & (new_n73_ | (new_n104_ & \a[5] ) | (~new_n104_ & ~\a[5] )) & (~new_n73_ | (new_n104_ ^ \a[5] ))) | (~\a[2]  & (new_n73_ ^ (new_n104_ ^ \a[5] ))))) | (\a[2]  & ((new_n72_ & \a[5] ) | (~new_n72_ & ~\a[5] ) | ((~new_n104_ | ~\a[5] ) & (new_n73_ | (new_n104_ & \a[5] ) | (~new_n104_ & ~\a[5] )))) & ((new_n72_ ^ \a[5] ) | (new_n104_ & \a[5] ) | (~new_n73_ & (~new_n104_ | ~\a[5] ) & (new_n104_ | \a[5] )))) | (~\a[2]  & ((~new_n72_ ^ \a[5] ) ^ ((new_n104_ & \a[5] ) | (~new_n73_ & (~new_n104_ | ~\a[5] ) & (new_n104_ | \a[5] ))))));
  assign new_n104_ = ~new_n48_ ^ new_n64_;
  assign new_n105_ = (new_n75_ ^ \a[5] ) ^ ((\a[5]  & (~new_n74_ | ((new_n54_ | ~new_n63_) & (new_n57_ | (~new_n54_ & new_n63_) | (new_n54_ & ~new_n63_)))) & (new_n74_ | (~new_n54_ & new_n63_) | (~new_n57_ & (new_n54_ | ~new_n63_) & (~new_n54_ | new_n63_)))) | ((~\a[5]  | (new_n74_ & ((~new_n54_ & new_n63_) | (~new_n57_ & (new_n54_ | ~new_n63_) & (~new_n54_ | new_n63_)))) | (~new_n74_ & (new_n54_ | ~new_n63_) & (new_n57_ | (~new_n54_ & new_n63_) | (new_n54_ & ~new_n63_)))) & (\a[5]  | (new_n74_ ^ ((~new_n54_ & new_n63_) | (~new_n57_ & (new_n54_ | ~new_n63_) & (~new_n54_ | new_n63_))))) & ((~new_n91_ & (new_n57_ | (~new_n54_ & new_n63_) | (new_n54_ & ~new_n63_)) & (~new_n57_ | (~new_n54_ ^ new_n63_))) | (~new_n76_ & (new_n91_ | (~new_n57_ & (new_n54_ | ~new_n63_) & (~new_n54_ | new_n63_)) | (new_n57_ & (new_n54_ ^ new_n63_))) & (~new_n91_ | (~new_n57_ ^ (~new_n54_ ^ new_n63_)))))));
  assign new_n106_ = (~\a[2]  | (new_n107_ & (new_n108_ | (~new_n76_ & new_n110_))) | (~new_n107_ & ~new_n108_ & (new_n76_ | ~new_n110_))) & (((~\a[2]  | (~new_n76_ & new_n110_) | (new_n76_ & ~new_n110_)) & (((~new_n111_ | ~\a[2] ) & ((new_n111_ & \a[2] ) | (~new_n111_ & ~\a[2] ) | ((~new_n112_ | ~\a[2] ) & (new_n113_ | (new_n112_ & \a[2] ) | (~new_n112_ & ~\a[2] ))))) | (\a[2]  & (new_n76_ | ~new_n110_) & (~new_n76_ | new_n110_)) | (~\a[2]  & (new_n76_ ^ new_n110_)))) | (\a[2]  & (~new_n107_ | (~new_n108_ & (new_n76_ | ~new_n110_))) & (new_n107_ | new_n108_ | (~new_n76_ & new_n110_))) | (~\a[2]  & (~new_n107_ ^ (new_n108_ | (~new_n76_ & new_n110_)))));
  assign new_n107_ = \a[5]  ^ ((~new_n52_ ^ new_n53_) ^ ((~new_n54_ & new_n63_) | (~new_n57_ & (new_n54_ | ~new_n63_) & (~new_n54_ | new_n63_))));
  assign new_n108_ = ~new_n91_ & (new_n57_ | ~new_n109_) & (~new_n57_ | new_n109_);
  assign new_n109_ = new_n63_ ^ (~\a[8]  ^ (new_n56_ & (~new_n33_ | ~new_n55_)));
  assign new_n110_ = ~new_n91_ ^ (~new_n57_ ^ new_n109_);
  assign new_n111_ = (~new_n77_ ^ new_n78_) ^ ((new_n79_ & ~new_n80_) | ((new_n79_ | ~new_n80_) & (~new_n79_ | new_n80_) & ((~new_n81_ & new_n90_) | (~new_n84_ & (new_n81_ | ~new_n90_) & (~new_n81_ | new_n90_)))));
  assign new_n112_ = (~new_n79_ ^ new_n80_) ^ ((~new_n81_ & new_n90_) | (~new_n84_ & (new_n81_ | ~new_n90_) & (~new_n81_ | new_n90_)));
  assign new_n113_ = (new_n115_ | (~new_n84_ & new_n114_) | (new_n84_ & ~new_n114_)) & ((~new_n115_ & (new_n84_ | ~new_n114_) & (~new_n84_ | new_n114_)) | (new_n115_ & (new_n84_ ^ new_n114_)) | ((new_n116_ | ~new_n117_) & ((~new_n116_ & new_n117_) | (new_n116_ & ~new_n117_) | (~new_n118_ & (new_n121_ | ~new_n127_)))));
  assign new_n114_ = new_n90_ ^ (~\a[5]  ^ (new_n83_ & (~new_n33_ | ~new_n82_)));
  assign new_n115_ = \a[2]  ^ (~\b[6]  | (((~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (new_n47_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))));
  assign new_n116_ = \a[2]  ^ (((new_n47_ ^ \b[6] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[5]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[6]  | \a[0]  | ~\a[1] ));
  assign new_n117_ = (new_n87_ | (~new_n88_ & new_n89_)) ^ (new_n86_ ^ (~\a[5]  ^ (new_n85_ & (~new_n36_ | ~new_n82_))));
  assign new_n118_ = (~\a[2]  ^ (new_n120_ & (~new_n30_ | ~new_n119_))) & (new_n88_ | ~new_n89_) & (~new_n88_ | new_n89_);
  assign new_n119_ = \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] );
  assign new_n120_ = (~\b[4]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[6]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[5]  | \a[0]  | ~\a[1] );
  assign new_n121_ = (~new_n123_ | (\a[2]  ^ (new_n122_ & (~new_n33_ | ~new_n119_)))) & ((new_n123_ & (~\a[2]  ^ (new_n122_ & (~new_n33_ | ~new_n119_)))) | (~new_n123_ & (~\a[2]  | ~new_n122_ | (new_n33_ & new_n119_)) & (\a[2]  | (new_n122_ & (~new_n33_ | ~new_n119_)))) | ((new_n124_ | ~new_n125_) & (~new_n126_ | (~new_n124_ & new_n125_) | (new_n124_ & ~new_n125_))));
  assign new_n122_ = (~\b[3]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[5]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[4]  | \a[0]  | ~\a[1] );
  assign new_n123_ = (~\a[5]  | ((~\b[0]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[5]  & (~\b[0]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] )))) ^ ((~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (\a[2]  ^ \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )) & (~\b[1]  | (\a[2]  ^ \a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[2]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n124_ = \a[2]  ^ ((~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )))) | ((~\b[3]  ^ \b[4] ) & (~\b[2]  | ~\b[3] ) & ((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[4]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[3]  | \a[0]  | ~\a[1] ));
  assign new_n125_ = ((\b[0]  & (~\a[2]  ^ \a[3] ) & (\a[3]  | \a[4] ) & (~\a[3]  | ~\a[4] )) | (\b[1]  & (~\a[2]  | ~\a[3] ) & (\a[2]  | \a[3] ) & (\a[4]  ^ ~\a[5] )) | ((~\a[2]  | ~\a[3] ) & (\a[2]  | \a[3] ) & (\a[4]  | \a[5] ) & (~\a[4]  | ~\a[5] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[5]  & \b[0]  & (~\a[2]  | ~\a[3] ) & (\a[2]  | \a[3] ));
  assign new_n126_ = ((\b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] )) | (\a[2]  & (~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] ) & (((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))) | (~\a[2]  & ((\b[1]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[3]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[2]  & ~\a[0]  & \a[1] ) | (((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )) & ((\b[2]  ^ \b[3] ) | (\b[1]  & (\b[0]  | \b[2] ))) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] ))))) & ((\b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (~\a[2]  ^ ((~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] ) & (((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))))) | (\a[2]  & (~\b[1]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[0]  | \a[0]  | ~\a[1] ) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\a[0]  | ~\b[0] ) & (~\b[2]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[1]  | \a[0]  | ~\a[1] ) & (~\b[0]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & ((\b[2]  ^ (\b[0]  | ~\b[1] )) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))));
  assign new_n127_ = (~\a[2]  ^ (new_n120_ & (~new_n30_ | ~new_n119_))) ^ (~new_n88_ ^ new_n89_);
  assign new_n128_ = ((\a[2]  & (new_n73_ | (new_n104_ & \a[5] ) | (~new_n104_ & ~\a[5] )) & (~new_n73_ | (new_n104_ ^ \a[5] ))) | (((new_n105_ & \a[2] ) | (~new_n106_ & (~new_n105_ | ~\a[2] ) & (new_n105_ | \a[2] ))) & (~\a[2]  | (~new_n73_ & (~new_n104_ | ~\a[5] ) & (new_n104_ | \a[5] )) | (new_n73_ & (~new_n104_ ^ \a[5] ))) & (\a[2]  | (~new_n73_ ^ (new_n104_ ^ \a[5] ))))) ^ (\a[2]  ^ ((new_n72_ ^ \a[5] ) ^ ((new_n104_ & \a[5] ) | (~new_n73_ & (~new_n104_ | ~\a[5] ) & (new_n104_ | \a[5] )))));
  assign new_n129_ = ((~\a[2]  ^ (~new_n73_ ^ new_n130_)) ^ ((new_n105_ & \a[2] ) | ((~new_n105_ | ~\a[2] ) & (new_n105_ | \a[2] ) & ((new_n131_ & \a[2] ) | ((~new_n131_ | ~\a[2] ) & (new_n131_ | \a[2] ) & ((new_n132_ & \a[2] ) | (~new_n133_ & (~new_n132_ | ~\a[2] ) & (new_n132_ | \a[2] )))))))) & ((new_n105_ ^ \a[2] ) | (new_n131_ & \a[2] ) | ((~new_n131_ | ~\a[2] ) & (new_n131_ | \a[2] ) & ((new_n132_ & \a[2] ) | (~new_n133_ & (~new_n132_ | ~\a[2] ) & (new_n132_ | \a[2] ))))) & ((new_n105_ & \a[2] ) | (~new_n105_ & ~\a[2] ) | ((~new_n131_ | ~\a[2] ) & ((new_n131_ & \a[2] ) | (~new_n131_ & ~\a[2] ) | ((~new_n132_ | ~\a[2] ) & (new_n133_ | (new_n132_ & \a[2] ) | (~new_n132_ & ~\a[2] )))))) & ((~new_n131_ ^ \a[2] ) ^ ((new_n132_ & \a[2] ) | (~new_n133_ & (~new_n132_ | ~\a[2] ) & (new_n132_ | \a[2] )))) & new_n135_ & (new_n133_ ^ (new_n132_ ^ \a[2] ));
  assign new_n130_ = \a[5]  ^ (~new_n48_ ^ new_n64_);
  assign new_n131_ = new_n107_ ^ (new_n108_ | (~new_n76_ & new_n110_));
  assign new_n132_ = ~new_n76_ ^ new_n110_;
  assign new_n133_ = (~new_n111_ | ~\a[2] ) & (~new_n134_ | ((~new_n112_ | ~\a[2] ) & (new_n113_ | (new_n112_ & \a[2] ) | (~new_n112_ & ~\a[2] ))));
  assign new_n134_ = \a[2]  ^ ((~new_n77_ ^ new_n78_) ^ ((new_n79_ & ~new_n80_) | ((new_n79_ | ~new_n80_) & (~new_n79_ | new_n80_) & ((~new_n81_ & new_n90_) | (~new_n84_ & (new_n81_ | ~new_n90_) & (~new_n81_ | new_n90_))))));
  assign new_n135_ = (new_n134_ | (new_n112_ & \a[2] ) | (~new_n113_ & (~new_n112_ | ~\a[2] ) & (new_n112_ | \a[2] ))) & (~new_n134_ | ((~new_n112_ | ~\a[2] ) & (new_n113_ | (new_n112_ & \a[2] ) | (~new_n112_ & ~\a[2] )))) & (~new_n113_ | (new_n112_ ^ \a[2] )) & (new_n113_ | (new_n112_ & \a[2] ) | (~new_n112_ & ~\a[2] )) & (~new_n136_ | new_n137_) & new_n138_ & (new_n136_ | ~new_n137_);
  assign new_n136_ = (new_n116_ | ~new_n117_) & ((~new_n118_ & (new_n121_ | ~new_n127_)) | (~new_n116_ & new_n117_) | (new_n116_ & ~new_n117_));
  assign new_n137_ = ~new_n115_ ^ (~new_n84_ ^ new_n114_);
  assign new_n138_ = ((~new_n118_ & (new_n121_ | ~new_n127_)) ^ (~new_n116_ ^ new_n117_)) & (new_n121_ ^ new_n127_) & ~new_n139_ & ~new_n140_ & new_n141_;
  assign new_n139_ = (new_n123_ ^ (~\a[2]  ^ (new_n122_ & (~new_n33_ | ~new_n119_)))) ^ ((~new_n124_ & new_n125_) | (new_n126_ & (new_n124_ | ~new_n125_) & (~new_n124_ | new_n125_)));
  assign new_n140_ = new_n126_ ^ (~new_n124_ ^ new_n125_);
  assign new_n141_ = ~new_n144_ & ~new_n145_ & (new_n143_ | ~\a[2] ) & new_n147_ & (~new_n146_ | ~new_n142_ | \a[1]  | \a[2] );
  assign new_n142_ = ~\a[9]  & ~\a[10] ;
  assign new_n143_ = (~\b[2]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[1]  | \a[0]  | ~\a[1] ) & (~\b[0]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )));
  assign new_n144_ = (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) ^ (\a[2]  ^ ((~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] ) & (((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))));
  assign new_n145_ = (((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[1]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[0]  | \a[0]  | ~\a[1] )) ? ~\a[2]  : ((~\b[2]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[1]  | \a[0]  | ~\a[1] ) & (~\b[0]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n146_ = ~\a[5]  & ~\a[6]  & ~\a[11]  & ~\a[12]  & ~\a[3]  & ~\a[4]  & ~\a[7]  & ~\a[8] ;
  assign new_n147_ = \a[0]  & \b[0]  & (\b[5]  | \b[6]  | \b[2]  | \b[3]  | \b[1]  | \b[4] );
endmodule


