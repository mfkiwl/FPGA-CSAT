// Benchmark "multiplier_999999000001_sat" written by ABC on Fri Nov 11 19:05:46 2022

module multiplier_999999000001_sat ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \b[0] , \b[1] ,
    \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] ,
    sat  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] ;
  output sat;
  wire new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_,
    new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_,
    new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_, new_n83_,
    new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_,
    new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_,
    new_n98_, new_n99_, new_n100_, new_n101_, new_n102_, new_n103_,
    new_n104_, new_n105_, new_n106_, new_n107_, new_n108_, new_n109_,
    new_n110_, new_n111_, new_n112_, new_n113_, new_n114_, new_n115_,
    new_n116_, new_n117_, new_n118_, new_n119_, new_n120_, new_n121_,
    new_n122_, new_n123_, new_n124_, new_n125_, new_n126_, new_n127_,
    new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_,
    new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_,
    new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_,
    new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_,
    new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_,
    new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_,
    new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_,
    new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_,
    new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_,
    new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_,
    new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_,
    new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_,
    new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_,
    new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_,
    new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_,
    new_n1166_, new_n1167_;
  assign sat = ~new_n1098_ & new_n1099_ & ((~new_n63_ ^ ~new_n906_) ^ (~new_n1010_ ^ (~new_n1167_ ^ (\a[5]  ^ ~\a[8] ))));
  assign new_n63_ = ~new_n900_ ^ (~new_n64_ ^ new_n905_);
  assign new_n64_ = (~\a[8]  | (((new_n894_ & \a[11] ) | ((~new_n894_ | ~\a[11] ) & (new_n894_ | \a[11] ) & ((new_n897_ & \a[11] ) | (~new_n898_ & (~new_n897_ | ~\a[11] ) & (new_n897_ | \a[11] ))))) & (~\a[11]  | (new_n65_ & ~new_n899_) | (~new_n65_ & new_n899_)) & (\a[11]  | (new_n65_ ^ ~new_n899_))) | ((~new_n894_ | ~\a[11] ) & ((new_n894_ & \a[11] ) | (~new_n894_ & ~\a[11] ) | ((~new_n897_ | ~\a[11] ) & (new_n898_ | (new_n897_ & \a[11] ) | (~new_n897_ & ~\a[11] )))) & (~\a[11]  ^ (new_n65_ ^ ~new_n899_)))) & (((~\a[8]  | ((~new_n894_ | ~\a[11] ) & (new_n894_ | \a[11] ) & ((new_n897_ & \a[11] ) | (~new_n898_ & (~new_n897_ | ~\a[11] ) & (new_n897_ | \a[11] )))) | ((~new_n894_ ^ \a[11] ) & (~new_n897_ | ~\a[11] ) & (new_n898_ | (new_n897_ & \a[11] ) | (~new_n897_ & ~\a[11] )))) & ((\a[8]  & ((new_n894_ & \a[11] ) | (~new_n894_ & ~\a[11] ) | ((~new_n897_ | ~\a[11] ) & (new_n898_ | (new_n897_ & \a[11] ) | (~new_n897_ & ~\a[11] )))) & ((new_n894_ ^ \a[11] ) | (new_n897_ & \a[11] ) | (~new_n898_ & (~new_n897_ | ~\a[11] ) & (new_n897_ | \a[11] )))) | (~\a[8]  & ((~new_n894_ ^ \a[11] ) ^ ((new_n897_ & \a[11] ) | (~new_n898_ & (~new_n897_ | ~\a[11] ) & (new_n897_ | \a[11] ))))) | ((~\a[8]  | (~new_n898_ & (~new_n897_ | ~\a[11] ) & (new_n897_ | \a[11] )) | (new_n898_ & (~new_n897_ ^ \a[11] ))) & (new_n640_ | (\a[8]  & (new_n898_ | (new_n897_ & \a[11] ) | (~new_n897_ & ~\a[11] )) & (~new_n898_ | (new_n897_ ^ \a[11] ))) | (~\a[8]  & (new_n898_ ^ (new_n897_ ^ \a[11] ))))))) | (\a[8]  & (((~new_n894_ | ~\a[11] ) & ((new_n894_ & \a[11] ) | (~new_n894_ & ~\a[11] ) | ((~new_n897_ | ~\a[11] ) & (new_n898_ | (new_n897_ & \a[11] ) | (~new_n897_ & ~\a[11] ))))) | (\a[11]  & (~new_n65_ | new_n899_) & (new_n65_ | ~new_n899_)) | (~\a[11]  & (~new_n65_ ^ ~new_n899_))) & ((new_n894_ & \a[11] ) | ((~new_n894_ | ~\a[11] ) & (new_n894_ | \a[11] ) & ((new_n897_ & \a[11] ) | (~new_n898_ & (~new_n897_ | ~\a[11] ) & (new_n897_ | \a[11] )))) | (\a[11]  ^ (new_n65_ ^ ~new_n899_)))) | (~\a[8]  & (((~new_n894_ | ~\a[11] ) & ((new_n894_ & \a[11] ) | (~new_n894_ & ~\a[11] ) | ((~new_n897_ | ~\a[11] ) & (new_n898_ | (new_n897_ & \a[11] ) | (~new_n897_ & ~\a[11] ))))) ^ (\a[11]  ^ (new_n65_ ^ ~new_n899_)))));
  assign new_n65_ = \a[14]  ^ (new_n66_ ^ ~new_n561_);
  assign new_n66_ = \a[17]  ^ (((new_n560_ & \a[20] ) | (~new_n67_ & (~new_n560_ | ~\a[20] ) & (new_n560_ | \a[20] ))) ^ (~new_n544_ ^ ~\a[20] ));
  assign new_n67_ = (~new_n531_ | ~\a[20] ) & (new_n68_ | (new_n531_ & \a[20] ) | (~new_n531_ & ~\a[20] ));
  assign new_n68_ = (~new_n494_ | ~\a[20] ) & ((new_n494_ & \a[20] ) | (~new_n494_ & ~\a[20] ) | ((~\a[20]  | ((new_n508_ | \a[23] ) & (~new_n508_ | ~\a[23] ) & ((new_n495_ & \a[23] ) | (~new_n507_ & (~new_n495_ | ~\a[23] ) & (new_n495_ | \a[23] )))) | ((new_n508_ ^ ~\a[23] ) & (~new_n495_ | ~\a[23] ) & (new_n507_ | (new_n495_ & \a[23] ) | (~new_n495_ & ~\a[23] )))) & (((~\a[20]  | (~new_n507_ & (~new_n495_ | ~\a[23] ) & (new_n495_ | \a[23] )) | (new_n507_ & (~new_n495_ ^ \a[23] ))) & (new_n69_ | (\a[20]  & (new_n507_ | (new_n495_ & \a[23] ) | (~new_n495_ & ~\a[23] )) & (~new_n507_ | (new_n495_ ^ \a[23] ))) | (~\a[20]  & (new_n507_ ^ (new_n495_ ^ \a[23] ))))) | (\a[20]  & ((~new_n508_ & ~\a[23] ) | (new_n508_ & \a[23] ) | ((~new_n495_ | ~\a[23] ) & (new_n507_ | (new_n495_ & \a[23] ) | (~new_n495_ & ~\a[23] )))) & ((~new_n508_ ^ ~\a[23] ) | (new_n495_ & \a[23] ) | (~new_n507_ & (~new_n495_ | ~\a[23] ) & (new_n495_ | \a[23] )))) | (~\a[20]  & ((new_n508_ ^ ~\a[23] ) ^ ((new_n495_ & \a[23] ) | (~new_n507_ & (~new_n495_ | ~\a[23] ) & (new_n495_ | \a[23] ))))))));
  assign new_n69_ = (~new_n344_ | ~\a[20] ) & (((~\a[20]  | ((~new_n70_ | ~\a[23] ) & (new_n70_ | \a[23] ) & ((new_n361_ & \a[23] ) | ((~new_n361_ | ~\a[23] ) & (new_n361_ | \a[23] ) & ((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )))))) | ((~new_n70_ ^ \a[23] ) & (~new_n361_ | ~\a[23] ) & ((new_n361_ & \a[23] ) | (~new_n361_ & ~\a[23] ) | ((~new_n362_ | ~\a[23] ) & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )))))) & (((~\a[20]  | ((~new_n361_ | ~\a[23] ) & (new_n361_ | \a[23] ) & ((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )))) | ((~new_n361_ ^ \a[23] ) & (~new_n362_ | ~\a[23] ) & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )))) & ((\a[20]  & ((new_n361_ & \a[23] ) | (~new_n361_ & ~\a[23] ) | ((~new_n362_ | ~\a[23] ) & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )))) & ((new_n361_ ^ \a[23] ) | (new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )))) | (~\a[20]  & ((~new_n361_ ^ \a[23] ) ^ ((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] ))))) | ((~\a[20]  | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )) | (new_n363_ & (~new_n362_ ^ \a[23] ))) & (new_n429_ | (\a[20]  & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )) & (~new_n363_ | (new_n362_ ^ \a[23] ))) | (~\a[20]  & (new_n363_ ^ (new_n362_ ^ \a[23] ))))))) | (\a[20]  & ((new_n70_ & \a[23] ) | (~new_n70_ & ~\a[23] ) | ((~new_n361_ | ~\a[23] ) & ((new_n361_ & \a[23] ) | (~new_n361_ & ~\a[23] ) | ((~new_n362_ | ~\a[23] ) & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )))))) & ((new_n70_ ^ \a[23] ) | (new_n361_ & \a[23] ) | ((~new_n361_ | ~\a[23] ) & (new_n361_ | \a[23] ) & ((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )))))) | (~\a[20]  & ((~new_n70_ ^ \a[23] ) ^ ((new_n361_ & \a[23] ) | ((~new_n361_ | ~\a[23] ) & (new_n361_ | \a[23] ) & ((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] ))))))))) | (new_n344_ & \a[20] ) | (~new_n344_ & ~\a[20] ));
  assign new_n70_ = new_n71_ ^ ~new_n330_;
  assign new_n71_ = (~new_n72_ | ~\a[26] ) & (((~new_n267_ | ~\a[26] ) & ((new_n267_ & \a[26] ) | (~new_n267_ & ~\a[26] ) | ((~\a[26]  | (~new_n202_ & new_n329_) | (new_n202_ & ~new_n329_)) & (new_n268_ | (\a[26]  & (new_n202_ | ~new_n329_) & (~new_n202_ | new_n329_)) | (~\a[26]  & (new_n202_ ^ new_n329_)))))) | (new_n72_ & \a[26] ) | (~new_n72_ & ~\a[26] ));
  assign new_n72_ = new_n256_ ^ (new_n73_ | (new_n255_ & ((~new_n266_ & (new_n145_ | ~new_n188_) & (~new_n145_ | new_n188_)) | (~new_n202_ & (new_n266_ | (~new_n145_ & new_n188_) | (new_n145_ & ~new_n188_)) & (~new_n266_ | (~new_n145_ ^ new_n188_))))));
  assign new_n73_ = ~new_n200_ & (~new_n189_ | (~new_n74_ & (new_n145_ | ~new_n188_))) & (new_n189_ | new_n74_ | (~new_n145_ & new_n188_));
  assign new_n74_ = ~new_n143_ & (~new_n75_ | new_n136_) & (new_n75_ | ~new_n136_);
  assign new_n75_ = (~new_n76_ | new_n132_) & ((new_n76_ & ~new_n132_) | (~new_n76_ & new_n132_) | (~new_n105_ & (~new_n130_ | ((new_n134_ | (~new_n131_ & new_n85_) | (new_n131_ & ~new_n85_)) & (new_n108_ | (~new_n134_ & (new_n131_ | ~new_n85_) & (~new_n131_ | new_n85_)) | (new_n134_ & (new_n131_ ^ new_n85_)))))));
  assign new_n76_ = new_n77_ ^ (new_n103_ | (new_n82_ & (new_n84_ | new_n104_)));
  assign new_n77_ = ~new_n78_ ^ (\a[38]  & ~\b[7] );
  assign new_n78_ = new_n81_ & (~new_n80_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))))));
  assign new_n79_ = (~\b[6]  | ~\b[7] ) & (((~\b[5]  | ~\b[6] ) & ((\b[5]  & \b[6] ) | (~\b[5]  & ~\b[6] ) | ((~\b[4]  | ~\b[5] ) & ((\b[4]  & \b[5] ) | (~\b[4]  & ~\b[5] ) | ((~\b[3]  | ~\b[4] ) & ((\b[3]  & \b[4] ) | (~\b[3]  & ~\b[4] ) | ((~\b[2]  | ~\b[3] ) & ((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] ))))))))) | (\b[6]  & \b[7] ) | (~\b[6]  & ~\b[7] ));
  assign new_n80_ = (\a[35]  | \a[36] ) & (~\a[35]  | ~\a[36] ) & (~\a[37]  | ~\a[38] ) & (\a[37]  | \a[38] );
  assign new_n81_ = (~\b[8]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (~\a[35]  ^ ~\a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[9]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[10]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] ));
  assign new_n82_ = ~new_n83_ ^ (\a[38]  & ~\b[6] );
  assign new_n83_ = (((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))) | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] )) & (~\b[7]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (\a[35]  ^ \a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[8]  | (\a[35]  ^ \a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[9]  | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  ^ \a[38] ));
  assign new_n84_ = new_n85_ & (new_n102_ | (new_n87_ & (new_n101_ | (new_n90_ & (new_n100_ | (new_n93_ & ~new_n96_))))));
  assign new_n85_ = (\a[38]  & ~\b[5] ) ^ (~new_n86_ | (new_n80_ & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )) & (~new_n79_ | (\b[7]  ^ \b[8] ))));
  assign new_n86_ = (~\b[6]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (~\a[35]  ^ ~\a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[7]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[8]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] ));
  assign new_n87_ = (\a[38]  & ~\b[4] ) ^ (~new_n89_ | (new_n80_ & new_n88_));
  assign new_n88_ = ((\b[5]  & \b[6] ) | ((~\b[5]  | ~\b[6] ) & (\b[5]  | \b[6] ) & ((\b[4]  & \b[5] ) | ((~\b[4]  | ~\b[5] ) & (\b[4]  | \b[5] ) & ((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))))))) ^ (\b[6]  ^ \b[7] );
  assign new_n89_ = (~\b[5]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (~\a[35]  ^ ~\a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[6]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[7]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] ));
  assign new_n90_ = (\a[38]  & ~\b[3] ) ^ (~new_n92_ | (new_n80_ & new_n91_));
  assign new_n91_ = (\b[5]  ^ \b[6] ) ^ ((\b[4]  & \b[5] ) | ((~\b[4]  | ~\b[5] ) & (\b[4]  | \b[5] ) & ((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )))))));
  assign new_n92_ = (~\b[4]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (~\a[35]  ^ ~\a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[5]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[6]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] ));
  assign new_n93_ = (\a[38]  & ~\b[2] ) ^ (~new_n95_ | (new_n80_ & new_n94_));
  assign new_n94_ = (\b[4]  ^ \b[5] ) ^ ((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )))));
  assign new_n95_ = (~\b[3]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (~\a[35]  ^ ~\a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[4]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[5]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] ));
  assign new_n96_ = (new_n97_ | (\a[38]  & ~\b[1]  & (~new_n99_ | (new_n80_ & new_n98_))) | ((~\a[38]  | \b[1] ) & new_n99_ & (~new_n80_ | ~new_n98_))) & (~\a[38]  | ~\b[1]  | ~new_n99_ | (new_n80_ & new_n98_));
  assign new_n97_ = (~\a[38]  | ~\b[0]  | (\b[0]  & (\a[35]  ^ ~\a[36] ) & (~\a[36]  | ~\a[37] ) & (\a[36]  | \a[37] )) | (\b[1]  & (\a[35]  | \a[36] ) & (~\a[35]  | ~\a[36] ) & (~\a[37]  ^ \a[38] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & (\a[35]  | \a[36] ) & (~\a[35]  | ~\a[36] ) & (~\a[37]  | ~\a[38] ) & (\a[37]  | \a[38] )) | (\b[0]  & (\a[35]  | \a[36] ) & (~\a[35]  | ~\a[36] )) | (\b[0]  & (~\a[37]  | ~\a[38] ) & (\a[37]  | \a[38] ) & (\a[35]  ^ ~\a[36] ) & (~\a[36]  ^ \a[37] )) | (\b[1]  & (\a[35]  ^ ~\a[36] ) & (~\a[36]  | ~\a[37] ) & (\a[36]  | \a[37] )) | (\b[2]  & (\a[35]  | \a[36] ) & (~\a[35]  | ~\a[36] ) & (~\a[37]  ^ \a[38] )) | ((\a[35]  | \a[36] ) & (~\a[35]  | ~\a[36] ) & (~\a[37]  | ~\a[38] ) & (\a[37]  | \a[38] ) & (~\b[2]  ^ (\b[0]  | ~\b[1] )))) & ((\a[38]  ^ (((~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (~\a[35]  ^ ~\a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[2]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[3]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] )))) | (\a[38]  & \b[0]  & (~\b[0]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[1]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] )) & (~\b[0]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] )) & (~\b[0]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (~\a[35]  ^ ~\a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[1]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[2]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] )) & ((~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))) | ((~\a[38]  | ~\b[0] ) & ((\b[0]  & (\a[35]  ^ ~\a[36] ) & (~\a[36]  | ~\a[37] ) & (\a[36]  | \a[37] )) | (\b[1]  & (\a[35]  | \a[36] ) & (~\a[35]  | ~\a[36] ) & (~\a[37]  ^ \a[38] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & (\a[35]  | \a[36] ) & (~\a[35]  | ~\a[36] ) & (~\a[37]  | ~\a[38] ) & (\a[37]  | \a[38] )) | ~\a[38]  | (\b[0]  & (\a[35]  | \a[36] ) & (~\a[35]  | ~\a[36] )) | (\b[0]  & (~\a[37]  | ~\a[38] ) & (\a[37]  | \a[38] ) & (\a[35]  ^ ~\a[36] ) & (~\a[36]  ^ \a[37] )) | (\b[1]  & (\a[35]  ^ ~\a[36] ) & (~\a[36]  | ~\a[37] ) & (\a[36]  | \a[37] )) | (\b[2]  & (\a[35]  | \a[36] ) & (~\a[35]  | ~\a[36] ) & (~\a[37]  ^ \a[38] )) | ((\a[35]  | \a[36] ) & (~\a[35]  | ~\a[36] ) & (~\a[37]  | ~\a[38] ) & (\a[37]  | \a[38] ) & (~\b[2]  ^ (\b[0]  | ~\b[1] ))))));
  assign new_n98_ = (\b[3]  ^ \b[4] ) ^ ((\b[2]  & \b[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )));
  assign new_n99_ = (~\b[2]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (~\a[35]  ^ ~\a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[3]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[4]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] ));
  assign new_n100_ = \a[38]  & \b[2]  & new_n95_ & (~new_n80_ | ~new_n94_);
  assign new_n101_ = \a[38]  & \b[3]  & new_n92_ & (~new_n80_ | ~new_n91_);
  assign new_n102_ = \a[38]  & \b[4]  & new_n89_ & (~new_n80_ | ~new_n88_);
  assign new_n103_ = new_n83_ & \a[38]  & \b[6] ;
  assign new_n104_ = \a[38]  & \b[5]  & new_n86_ & (~new_n80_ | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n79_ & (~\b[7]  ^ \b[8] )));
  assign new_n105_ = ~new_n106_ & (~new_n82_ | (~new_n84_ & ~new_n104_)) & (new_n82_ | new_n84_ | new_n104_);
  assign new_n106_ = \a[35]  ^ ((~new_n107_ | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & (~\b[11]  | (\a[32]  ^ \a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[12]  | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[10]  | (\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )));
  assign new_n107_ = (\b[11]  ^ \b[12] ) ^ ((\b[10]  & \b[11] ) | ((~\b[10]  | ~\b[11] ) & (\b[10]  | \b[11] ) & ((\b[9]  & \b[10] ) | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | (((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))) & (~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] )))))));
  assign new_n108_ = (~new_n109_ | new_n127_) & ((~new_n110_ & (~new_n126_ | ((new_n129_ | (~new_n93_ & new_n96_) | (new_n93_ & ~new_n96_)) & (new_n112_ | (~new_n129_ & (new_n93_ | ~new_n96_) & (~new_n93_ | new_n96_)) | (new_n129_ & (new_n93_ ^ new_n96_)))))) | (new_n109_ & ~new_n127_) | (~new_n109_ & new_n127_));
  assign new_n109_ = new_n87_ ^ (new_n101_ | (new_n90_ & (new_n100_ | (new_n93_ & ~new_n96_))));
  assign new_n110_ = ~new_n111_ & (~new_n90_ | (~new_n100_ & (~new_n93_ | new_n96_))) & (new_n90_ | new_n100_ | (new_n93_ & ~new_n96_));
  assign new_n111_ = \a[35]  ^ ((((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))) | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & (~\b[8]  | (\a[32]  ^ \a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[9]  | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[7]  | (\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )));
  assign new_n112_ = (~new_n113_ | new_n114_) & ((new_n113_ & ~new_n114_) | (~new_n113_ & new_n114_) | ((new_n115_ | ~new_n124_) & (((new_n116_ | ~new_n125_) & (new_n117_ | (~new_n116_ & new_n125_) | (new_n116_ & ~new_n125_))) | (~new_n115_ & new_n124_) | (new_n115_ & ~new_n124_))));
  assign new_n113_ = ~new_n97_ ^ ((\a[38]  & ~\b[1] ) ^ (~new_n99_ | (new_n80_ & new_n98_)));
  assign new_n114_ = \a[35]  ^ ((~new_n88_ | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & (~\b[6]  | (\a[32]  ^ \a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[7]  | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[5]  | (\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )));
  assign new_n115_ = \a[35]  ^ ((~new_n91_ | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & (~\b[5]  | (\a[32]  ^ \a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[6]  | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[4]  | (\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )));
  assign new_n116_ = \a[35]  ^ ((~new_n94_ | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & (~\b[4]  | (\a[32]  ^ \a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[5]  | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[3]  | (\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )));
  assign new_n117_ = (~new_n120_ | (\a[35]  ^ (new_n119_ & (~new_n118_ | ~new_n98_)))) & ((~new_n121_ & (new_n122_ | ~new_n123_)) | (new_n120_ & (~\a[35]  ^ (new_n119_ & (~new_n118_ | ~new_n98_)))) | (~new_n120_ & (~\a[35]  | ~new_n119_ | (new_n118_ & new_n98_)) & (\a[35]  | (new_n119_ & (~new_n118_ | ~new_n98_)))));
  assign new_n118_ = (\a[32]  | \a[33] ) & (~\a[32]  | ~\a[33] ) & (~\a[34]  | ~\a[35] ) & (\a[34]  | \a[35] );
  assign new_n119_ = (~\b[3]  | (~\a[32]  ^ ~\a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[4]  | (~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[2]  | (\a[33]  ^ \a[34] ) | (~\a[32]  ^ ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] ));
  assign new_n120_ = ((\b[0]  & (\a[35]  ^ ~\a[36] ) & (~\a[36]  | ~\a[37] ) & (\a[36]  | \a[37] )) | (\b[1]  & (\a[35]  | \a[36] ) & (~\a[35]  | ~\a[36] ) & (~\a[37]  ^ \a[38] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & (\a[35]  | \a[36] ) & (~\a[35]  | ~\a[36] ) & (~\a[37]  | ~\a[38] ) & (\a[37]  | \a[38] ))) ^ ((\a[35]  | \a[36] ) & (~\a[35]  | ~\a[36] ) & \a[38]  & \b[0] );
  assign new_n121_ = \b[0]  & (~\a[35]  | ~\a[36] ) & (\a[35]  | \a[36] ) & (~\b[0]  | (~\a[32]  ^ ~\a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[1]  | (~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  ^ \a[35] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & \a[35]  & (~\b[0]  | (~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] )) & (~\b[0]  | (\a[33]  ^ \a[34] ) | (~\a[32]  ^ ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & (~\b[1]  | (~\a[32]  ^ ~\a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[2]  | (~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  ^ \a[35] )) & ((~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )));
  assign new_n122_ = \a[35]  ^ (((~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (~\a[32]  ^ ~\a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[3]  | (~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[1]  | (\a[33]  ^ \a[34] ) | (~\a[32]  ^ ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )));
  assign new_n123_ = (\b[0]  & (~\a[35]  | ~\a[36] ) & (\a[35]  | \a[36] )) ^ ((~\b[0]  | (~\a[32]  ^ ~\a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[1]  | (~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  ^ \a[35] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & \a[35]  & (~\b[0]  | (~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] )) & (~\b[0]  | (\a[33]  ^ \a[34] ) | (~\a[32]  ^ ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & (~\b[1]  | (~\a[32]  ^ ~\a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[2]  | (~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  ^ \a[35] )) & ((~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n124_ = (~\a[38]  ^ (((~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (~\a[35]  ^ ~\a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[2]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[3]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] )))) ^ ((\a[38]  & \b[0] ) ^ ((~\b[0]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[1]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] )) & \a[38]  & (~\b[0]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] )) & (~\b[0]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (~\a[35]  ^ ~\a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[1]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[2]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] )) & ((~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))));
  assign new_n125_ = ((~\b[0]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (~\a[35]  ^ ~\a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[1]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[2]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] )) & ((~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))) ^ (~\a[38]  | ((~\b[0]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[1]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] )) & \a[38]  & (~\b[0]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ))));
  assign new_n126_ = ~new_n111_ ^ (new_n90_ ^ (new_n100_ | (new_n93_ & ~new_n96_)));
  assign new_n127_ = \a[35]  ^ (new_n128_ & (~new_n118_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n128_ = (~\b[9]  | (~\a[32]  ^ ~\a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[10]  | (~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[8]  | (\a[33]  ^ \a[34] ) | (~\a[32]  ^ ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] ));
  assign new_n129_ = \a[35]  ^ ((~\b[7]  | (\a[32]  ^ \a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[8]  | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[6]  | (\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & ((\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n79_ & (~\b[7]  ^ \b[8] ))));
  assign new_n130_ = ~new_n106_ ^ (new_n82_ ^ (new_n84_ | new_n104_));
  assign new_n131_ = ~new_n102_ & (~new_n87_ | (~new_n101_ & (~new_n90_ | (~new_n100_ & (~new_n93_ | new_n96_)))));
  assign new_n132_ = \a[35]  ^ ((~new_n133_ | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & (~\b[12]  | (\a[32]  ^ \a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[13]  | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[11]  | (\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )));
  assign new_n133_ = (\b[12]  ^ \b[13] ) ^ ((\b[11]  & \b[12] ) | ((~\b[11]  | ~\b[12] ) & (\b[11]  | \b[12] ) & ((\b[10]  & \b[11] ) | ((~\b[10]  | ~\b[11] ) & (\b[10]  | \b[11] ) & ((\b[9]  & \b[10] ) | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | (((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))) & (~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] )))))))));
  assign new_n134_ = \a[35]  ^ ((~new_n135_ | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & (~\b[10]  | (\a[32]  ^ \a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[11]  | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[9]  | (\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )));
  assign new_n135_ = (\b[10]  ^ \b[11] ) ^ ((\b[9]  & \b[10] ) | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | (((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))) & (~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] )))));
  assign new_n136_ = ~new_n141_ ^ (new_n137_ ^ (new_n140_ | (new_n77_ & (new_n103_ | (new_n82_ & (new_n84_ | new_n104_))))));
  assign new_n137_ = ~new_n138_ ^ (\a[38]  & ~\b[8] );
  assign new_n138_ = new_n139_ & (~new_n80_ | ((~\b[10]  | ~\b[11] ) & (\b[10]  | \b[11] ) & ((\b[9]  & \b[10] ) | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))))) | ((~\b[10]  ^ \b[11] ) & (~\b[9]  | ~\b[10] ) & ((\b[9]  & \b[10] ) | (~\b[9]  & ~\b[10] ) | ((~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))))))));
  assign new_n139_ = (~\b[9]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (~\a[35]  ^ ~\a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[10]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[11]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] ));
  assign new_n140_ = new_n78_ & \a[38]  & \b[7] ;
  assign new_n141_ = \a[35]  ^ ((~\b[13]  | (\a[32]  ^ \a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[14]  | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[12]  | (\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & ((\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n142_ & (~\b[13]  ^ \b[14] ))));
  assign new_n142_ = (~\b[12]  | ~\b[13] ) & ((\b[12]  & \b[13] ) | (~\b[12]  & ~\b[13] ) | ((~\b[11]  | ~\b[12] ) & ((\b[11]  & \b[12] ) | (~\b[11]  & ~\b[12] ) | ((~\b[10]  | ~\b[11] ) & ((\b[10]  & \b[11] ) | (~\b[10]  & ~\b[11] ) | ((~\b[9]  | ~\b[10] ) & ((\b[9]  & \b[10] ) | (~\b[9]  & ~\b[10] ) | ((~\b[8]  | ~\b[9] ) & (((~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))) | (\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ))))))))));
  assign new_n143_ = \a[32]  ^ ((~new_n144_ | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & (~\b[16]  | (\a[29]  ^ \a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[17]  | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[15]  | (\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )));
  assign new_n144_ = (\b[16]  ^ \b[17] ) ^ ((\b[15]  & \b[16] ) | ((~\b[15]  | ~\b[16] ) & (\b[15]  | \b[16] ) & ((\b[14]  & \b[15] ) | (((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] ))) & (~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] )))));
  assign new_n145_ = (~new_n146_ | new_n185_) & ((~new_n150_ & (~new_n184_ | ((new_n187_ | (~new_n108_ & new_n148_) | (new_n108_ & ~new_n148_)) & (new_n152_ | (~new_n187_ & (new_n108_ | ~new_n148_) & (~new_n108_ | new_n148_)) | (new_n187_ & (new_n108_ ^ new_n148_)))))) | (new_n146_ & ~new_n185_) | (~new_n146_ & new_n185_));
  assign new_n146_ = new_n149_ ^ (new_n105_ | (new_n130_ & (new_n147_ | (~new_n108_ & new_n148_))));
  assign new_n147_ = ~new_n134_ & (new_n131_ | ~new_n85_) & (~new_n131_ | new_n85_);
  assign new_n148_ = ~new_n134_ ^ (~new_n131_ ^ new_n85_);
  assign new_n149_ = ~new_n132_ ^ (new_n77_ ^ (new_n103_ | (new_n82_ & (new_n84_ | new_n104_))));
  assign new_n150_ = ~new_n151_ & (~new_n130_ | (~new_n147_ & (new_n108_ | ~new_n148_))) & (new_n130_ | new_n147_ | (~new_n108_ & new_n148_));
  assign new_n151_ = \a[32]  ^ ((((~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] ) & ((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )))) | ((~\b[14]  ^ \b[15] ) & (~\b[13]  | ~\b[14] ) & (new_n142_ | (\b[13]  & \b[14] ) | (~\b[13]  & ~\b[14] ))) | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & (~\b[14]  | (\a[29]  ^ \a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[15]  | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[13]  | (\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )));
  assign new_n152_ = (~new_n153_ | new_n182_) & ((~new_n155_ & (~new_n180_ | ((new_n183_ | (~new_n112_ & new_n181_) | (new_n112_ & ~new_n181_)) & (new_n157_ | (~new_n183_ & (new_n112_ | ~new_n181_) & (~new_n112_ | new_n181_)) | (new_n183_ & (new_n112_ ^ new_n181_)))))) | (new_n153_ & ~new_n182_) | (~new_n153_ & new_n182_));
  assign new_n153_ = new_n154_ ^ (new_n110_ | (new_n126_ & ((~new_n129_ & (new_n93_ | ~new_n96_) & (~new_n93_ | new_n96_)) | (~new_n112_ & (new_n129_ | (~new_n93_ & new_n96_) | (new_n93_ & ~new_n96_)) & (~new_n129_ | (~new_n93_ ^ new_n96_))))));
  assign new_n154_ = ~new_n127_ ^ (new_n87_ ^ (new_n101_ | (new_n90_ & (new_n100_ | (new_n93_ & ~new_n96_)))));
  assign new_n155_ = ~new_n156_ & (~new_n126_ | ((new_n129_ | (~new_n93_ & new_n96_) | (new_n93_ & ~new_n96_)) & (new_n112_ | (~new_n129_ & (new_n93_ | ~new_n96_) & (~new_n93_ | new_n96_)) | (new_n129_ & (new_n93_ ^ new_n96_))))) & (new_n126_ | (~new_n129_ & (new_n93_ | ~new_n96_) & (~new_n93_ | new_n96_)) | (~new_n112_ & (new_n129_ | (~new_n93_ & new_n96_) | (new_n93_ & ~new_n96_)) & (~new_n129_ | (~new_n93_ ^ new_n96_))));
  assign new_n156_ = \a[32]  ^ ((~new_n107_ | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & (~\b[11]  | (\a[29]  ^ \a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[12]  | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[10]  | (\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )));
  assign new_n157_ = (~new_n159_ | new_n177_) & ((~new_n160_ & (~new_n176_ | ((new_n179_ | (new_n158_ & ~new_n117_) | (~new_n158_ & new_n117_)) & (new_n162_ | (~new_n179_ & (~new_n158_ | new_n117_) & (new_n158_ | ~new_n117_)) | (new_n179_ & (~new_n158_ ^ ~new_n117_)))))) | (new_n159_ & ~new_n177_) | (~new_n159_ & new_n177_));
  assign new_n158_ = new_n116_ ^ ~new_n125_;
  assign new_n159_ = (new_n113_ ^ ~new_n114_) ^ ((~new_n115_ & new_n124_) | (((~new_n116_ & new_n125_) | (~new_n117_ & (new_n116_ | ~new_n125_) & (~new_n116_ | new_n125_))) & (new_n115_ | ~new_n124_) & (~new_n115_ | new_n124_)));
  assign new_n160_ = ~new_n161_ & (((new_n116_ | ~new_n125_) & (new_n117_ | (~new_n116_ & new_n125_) | (new_n116_ & ~new_n125_))) | (~new_n115_ & new_n124_) | (new_n115_ & ~new_n124_)) & ((~new_n116_ & new_n125_) | (~new_n117_ & (new_n116_ | ~new_n125_) & (~new_n116_ | new_n125_)) | (~new_n115_ ^ new_n124_));
  assign new_n161_ = \a[32]  ^ ((((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))) | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & (~\b[8]  | (\a[29]  ^ \a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[9]  | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[7]  | (\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )));
  assign new_n162_ = (new_n163_ | ~new_n164_) & ((new_n163_ & ~new_n164_) | (~new_n163_ & new_n164_) | ((~new_n165_ | new_n166_) & (((new_n167_ | ~new_n175_) & (new_n168_ | (~new_n167_ & new_n175_) | (new_n167_ & ~new_n175_))) | (new_n165_ & ~new_n166_) | (~new_n165_ & new_n166_))));
  assign new_n163_ = \a[32]  ^ ((~new_n88_ | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & (~\b[6]  | (\a[29]  ^ \a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[7]  | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[5]  | (\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )));
  assign new_n164_ = (new_n121_ | (~new_n122_ & new_n123_)) ^ (new_n120_ ^ (~\a[35]  ^ (new_n119_ & (~new_n118_ | ~new_n98_))));
  assign new_n165_ = new_n122_ ^ ~new_n123_;
  assign new_n166_ = \a[32]  ^ ((~new_n91_ | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & (~\b[5]  | (\a[29]  ^ \a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[6]  | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[4]  | (\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )));
  assign new_n167_ = \a[32]  ^ ((~new_n94_ | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & (~\b[4]  | (\a[29]  ^ \a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[5]  | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[3]  | (\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )));
  assign new_n168_ = (~new_n171_ | (\a[32]  ^ (new_n170_ & (~new_n98_ | ~new_n169_)))) & ((~new_n172_ & (new_n173_ | ~new_n174_)) | (new_n171_ & (~\a[32]  ^ (new_n170_ & (~new_n98_ | ~new_n169_)))) | (~new_n171_ & (~\a[32]  | ~new_n170_ | (new_n98_ & new_n169_)) & (\a[32]  | (new_n170_ & (~new_n98_ | ~new_n169_)))));
  assign new_n169_ = (\a[29]  | \a[30] ) & (~\a[29]  | ~\a[30] ) & (~\a[31]  | ~\a[32] ) & (\a[31]  | \a[32] );
  assign new_n170_ = (~\b[3]  | (~\a[29]  ^ ~\a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[4]  | (~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[2]  | (\a[30]  ^ \a[31] ) | (~\a[29]  ^ ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] ));
  assign new_n171_ = ((\b[0]  & (\a[32]  ^ ~\a[33] ) & (~\a[33]  | ~\a[34] ) & (\a[33]  | \a[34] )) | (\b[1]  & (\a[32]  | \a[33] ) & (~\a[32]  | ~\a[33] ) & (~\a[34]  ^ \a[35] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & (\a[32]  | \a[33] ) & (~\a[32]  | ~\a[33] ) & (~\a[34]  | ~\a[35] ) & (\a[34]  | \a[35] ))) ^ (\a[35]  & \b[0]  & (\a[32]  | \a[33] ) & (~\a[32]  | ~\a[33] ));
  assign new_n172_ = \b[0]  & (~\a[32]  | ~\a[33] ) & (\a[32]  | \a[33] ) & (~\b[0]  | (~\a[29]  ^ ~\a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[1]  | (~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  ^ \a[32] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & \a[32]  & (~\b[0]  | (~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] )) & (~\b[0]  | (\a[30]  ^ \a[31] ) | (~\a[29]  ^ ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & (~\b[1]  | (~\a[29]  ^ ~\a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[2]  | (~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  ^ \a[32] )) & ((~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )));
  assign new_n173_ = \a[32]  ^ (((~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (~\a[29]  ^ ~\a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[3]  | (~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[1]  | (\a[30]  ^ \a[31] ) | (~\a[29]  ^ ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )));
  assign new_n174_ = (\b[0]  & (~\a[32]  | ~\a[33] ) & (\a[32]  | \a[33] )) ^ ((~\b[0]  | (~\a[29]  ^ ~\a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[1]  | (~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  ^ \a[32] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & \a[32]  & (~\b[0]  | (~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] )) & (~\b[0]  | (\a[30]  ^ \a[31] ) | (~\a[29]  ^ ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & (~\b[1]  | (~\a[29]  ^ ~\a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[2]  | (~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  ^ \a[32] )) & ((~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n175_ = (~\a[35]  | ((~\b[0]  | (~\a[32]  ^ ~\a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[1]  | (~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  ^ \a[35] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & \a[35]  & (~\b[0]  | (~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] )))) ^ ((~\b[1]  | (~\a[32]  ^ ~\a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[2]  | (~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  ^ \a[35] )) & ((~\a[32]  & ~\a[33] ) | (\a[32]  & \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (\a[33]  ^ \a[34] ) | (~\a[32]  ^ ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )));
  assign new_n176_ = ~new_n161_ ^ (((~new_n116_ & new_n125_) | (~new_n117_ & (new_n116_ | ~new_n125_) & (~new_n116_ | new_n125_))) ^ (~new_n115_ ^ new_n124_));
  assign new_n177_ = \a[32]  ^ (new_n178_ & (~new_n169_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n178_ = (~\b[9]  | (~\a[29]  ^ ~\a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[10]  | (~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[8]  | (\a[30]  ^ \a[31] ) | (~\a[29]  ^ ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] ));
  assign new_n179_ = \a[32]  ^ ((~\b[7]  | (\a[29]  ^ \a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[8]  | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[6]  | (\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & ((\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n79_ & (~\b[7]  ^ \b[8] ))));
  assign new_n180_ = ~new_n156_ ^ (new_n126_ ^ ((~new_n129_ & (new_n93_ | ~new_n96_) & (~new_n93_ | new_n96_)) | (~new_n112_ & (new_n129_ | (~new_n93_ & new_n96_) | (new_n93_ & ~new_n96_)) & (~new_n129_ | (~new_n93_ ^ new_n96_)))));
  assign new_n181_ = ~new_n129_ ^ (new_n93_ ^ ~new_n96_);
  assign new_n182_ = \a[32]  ^ ((~new_n133_ | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & (~\b[12]  | (\a[29]  ^ \a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[13]  | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[11]  | (\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )));
  assign new_n183_ = \a[32]  ^ ((~new_n135_ | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & (~\b[10]  | (\a[29]  ^ \a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[11]  | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[9]  | (\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )));
  assign new_n184_ = ~new_n151_ ^ (new_n130_ ^ (new_n147_ | (~new_n108_ & new_n148_)));
  assign new_n185_ = \a[32]  ^ ((~new_n186_ | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & (~\b[15]  | (\a[29]  ^ \a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[16]  | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[14]  | (\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )));
  assign new_n186_ = (\b[15]  ^ \b[16] ) ^ ((\b[14]  & \b[15] ) | (((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] ))) & (~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] )));
  assign new_n187_ = \a[32]  ^ ((~\b[13]  | (\a[29]  ^ \a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[14]  | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[12]  | (\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & ((\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n142_ & (~\b[13]  ^ \b[14] ))));
  assign new_n188_ = ~new_n143_ ^ (new_n75_ ^ ~new_n136_);
  assign new_n189_ = ~new_n198_ ^ (new_n191_ ^ (new_n190_ | new_n197_));
  assign new_n190_ = new_n136_ & ((new_n76_ & ~new_n132_) | ((new_n105_ | (new_n130_ & (new_n147_ | (~new_n108_ & new_n148_)))) & (~new_n76_ | new_n132_) & (new_n76_ | ~new_n132_)));
  assign new_n191_ = ~new_n196_ ^ (new_n192_ ^ ~new_n194_);
  assign new_n192_ = ~new_n193_ ^ (\a[38]  & ~\b[9] );
  assign new_n193_ = (~\b[10]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (\a[35]  ^ \a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[11]  | (\a[35]  ^ \a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[12]  | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  ^ \a[38] )) & (~new_n107_ | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ));
  assign new_n194_ = ~new_n195_ & (~new_n137_ | (~new_n140_ & (~new_n77_ | (~new_n103_ & (~new_n82_ | (~new_n84_ & ~new_n104_))))));
  assign new_n195_ = new_n138_ & \a[38]  & \b[8] ;
  assign new_n196_ = \a[35]  ^ ((((~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] ) & ((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )))) | ((~\b[14]  ^ \b[15] ) & (~\b[13]  | ~\b[14] ) & (new_n142_ | (\b[13]  & \b[14] ) | (~\b[13]  & ~\b[14] ))) | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & (~\b[14]  | (\a[32]  ^ \a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[15]  | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[13]  | (\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )));
  assign new_n197_ = ~new_n141_ & (~new_n137_ | (~new_n140_ & (~new_n77_ | (~new_n103_ & (~new_n82_ | (~new_n84_ & ~new_n104_)))))) & (new_n137_ | new_n140_ | (new_n77_ & (new_n103_ | (new_n82_ & (new_n84_ | new_n104_)))));
  assign new_n198_ = \a[32]  ^ ((~new_n199_ | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & (~\b[17]  | (\a[29]  ^ \a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[18]  | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[16]  | (\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )));
  assign new_n199_ = (\b[17]  ^ \b[18] ) ^ ((\b[16]  & \b[17] ) | ((~\b[16]  | ~\b[17] ) & (\b[16]  | \b[17] ) & ((\b[15]  & \b[16] ) | ((~\b[15]  | ~\b[16] ) & (\b[15]  | \b[16] ) & ((\b[14]  & \b[15] ) | (((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] ))) & (~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] )))))));
  assign new_n200_ = \a[29]  ^ (~\b[19]  | (((\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & (new_n201_ | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] ))));
  assign new_n201_ = (~\b[18]  | ~\b[19] ) & ((\b[18]  & \b[19] ) | (~\b[18]  & ~\b[19] ) | ((~\b[17]  | ~\b[18] ) & ((\b[17]  & \b[18] ) | (~\b[17]  & ~\b[18] ) | ((~\b[16]  | ~\b[17] ) & ((\b[16]  & \b[17] ) | (~\b[16]  & ~\b[17] ) | ((~\b[15]  | ~\b[16] ) & ((\b[15]  & \b[16] ) | (~\b[15]  & ~\b[16] ) | ((~\b[14]  | ~\b[15] ) & (((~\b[13]  | ~\b[14] ) & (new_n142_ | (\b[13]  & \b[14] ) | (~\b[13]  & ~\b[14] ))) | (\b[14]  & \b[15] ) | (~\b[14]  & ~\b[15] ))))))))));
  assign new_n202_ = (~new_n203_ | new_n252_) & ((~new_n207_ & (~new_n251_ | ((new_n254_ | (~new_n152_ & new_n205_) | (new_n152_ & ~new_n205_)) & (new_n209_ | (~new_n254_ & (new_n152_ | ~new_n205_) & (~new_n152_ | new_n205_)) | (new_n254_ & (new_n152_ ^ new_n205_)))))) | (new_n203_ & ~new_n252_) | (~new_n203_ & new_n252_));
  assign new_n203_ = new_n206_ ^ (new_n150_ | (new_n184_ & (new_n204_ | (~new_n152_ & new_n205_))));
  assign new_n204_ = ~new_n187_ & (~new_n108_ | new_n148_) & (new_n108_ | ~new_n148_);
  assign new_n205_ = ~new_n187_ ^ (new_n108_ ^ ~new_n148_);
  assign new_n206_ = ~new_n185_ ^ (new_n149_ ^ (new_n105_ | (new_n130_ & (new_n147_ | (~new_n108_ & new_n148_)))));
  assign new_n207_ = ~new_n208_ & (~new_n184_ | (~new_n204_ & (new_n152_ | ~new_n205_))) & (new_n184_ | new_n204_ | (~new_n152_ & new_n205_));
  assign new_n208_ = \a[29]  ^ ((~new_n199_ | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & (~\b[17]  | (\a[26]  ^ \a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[18]  | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[16]  | (\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )));
  assign new_n209_ = (~new_n210_ | new_n249_) & ((new_n210_ & ~new_n249_) | (~new_n210_ & new_n249_) | (~new_n214_ & (new_n214_ | new_n248_ | ((new_n250_ | (~new_n157_ & new_n212_) | (new_n157_ & ~new_n212_)) & (new_n216_ | (~new_n250_ & (new_n157_ | ~new_n212_) & (~new_n157_ | new_n212_)) | (new_n250_ & (new_n157_ ^ new_n212_)))))));
  assign new_n210_ = new_n213_ ^ (new_n155_ | (new_n180_ & (new_n211_ | (~new_n157_ & new_n212_))));
  assign new_n211_ = ~new_n183_ & (~new_n112_ | new_n181_) & (new_n112_ | ~new_n181_);
  assign new_n212_ = ~new_n183_ ^ (new_n112_ ^ ~new_n181_);
  assign new_n213_ = ~new_n182_ ^ (new_n154_ ^ (new_n110_ | (new_n126_ & ((~new_n129_ & (new_n93_ | ~new_n96_) & (~new_n93_ | new_n96_)) | (~new_n112_ & (new_n129_ | (~new_n93_ & new_n96_) | (new_n93_ & ~new_n96_)) & (~new_n129_ | (~new_n93_ ^ new_n96_)))))));
  assign new_n214_ = ~new_n215_ & (~new_n180_ | (~new_n211_ & (new_n157_ | ~new_n212_))) & (new_n180_ | new_n211_ | (~new_n157_ & new_n212_));
  assign new_n215_ = \a[29]  ^ ((((~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] ) & ((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )))) | ((~\b[14]  ^ \b[15] ) & (~\b[13]  | ~\b[14] ) & (new_n142_ | (\b[13]  & \b[14] ) | (~\b[13]  & ~\b[14] ))) | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & (~\b[14]  | (\a[26]  ^ \a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[15]  | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[13]  | (\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )));
  assign new_n216_ = (~new_n217_ | new_n246_) & ((new_n217_ & ~new_n246_) | (~new_n217_ & new_n246_) | (~new_n219_ & (~new_n221_ | ((new_n247_ | (~new_n162_ & new_n245_) | (new_n162_ & ~new_n245_)) & (new_n222_ | (~new_n247_ & (new_n162_ | ~new_n245_) & (~new_n162_ | new_n245_)) | (new_n247_ & (new_n162_ ^ new_n245_)))))));
  assign new_n217_ = new_n218_ ^ (new_n160_ | (new_n176_ & ((~new_n179_ & (new_n117_ | (~new_n116_ & new_n125_) | (new_n116_ & ~new_n125_)) & (~new_n117_ | (~new_n116_ ^ new_n125_))) | (~new_n162_ & (new_n179_ | (~new_n117_ & (new_n116_ | ~new_n125_) & (~new_n116_ | new_n125_)) | (new_n117_ & (new_n116_ ^ new_n125_))) & (~new_n179_ | (~new_n117_ ^ (~new_n116_ ^ new_n125_)))))));
  assign new_n218_ = ~new_n177_ ^ ((new_n113_ ^ ~new_n114_) ^ ((~new_n115_ & new_n124_) | (((~new_n116_ & new_n125_) | (~new_n117_ & (new_n116_ | ~new_n125_) & (~new_n116_ | new_n125_))) & (new_n115_ | ~new_n124_) & (~new_n115_ | new_n124_))));
  assign new_n219_ = ~new_n220_ & (~new_n176_ | ((new_n179_ | (~new_n117_ & (new_n116_ | ~new_n125_) & (~new_n116_ | new_n125_)) | (new_n117_ & (new_n116_ ^ new_n125_))) & (new_n162_ | (~new_n179_ & (new_n117_ | (~new_n116_ & new_n125_) | (new_n116_ & ~new_n125_)) & (~new_n117_ | (~new_n116_ ^ new_n125_))) | (new_n179_ & (new_n117_ ^ (~new_n116_ ^ new_n125_)))))) & (new_n176_ | (~new_n179_ & (new_n117_ | (~new_n116_ & new_n125_) | (new_n116_ & ~new_n125_)) & (~new_n117_ | (~new_n116_ ^ new_n125_))) | (~new_n162_ & (new_n179_ | (~new_n117_ & (new_n116_ | ~new_n125_) & (~new_n116_ | new_n125_)) | (new_n117_ & (new_n116_ ^ new_n125_))) & (~new_n179_ | (~new_n117_ ^ (~new_n116_ ^ new_n125_)))));
  assign new_n220_ = \a[29]  ^ ((~new_n107_ | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & (~\b[11]  | (\a[26]  ^ \a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[12]  | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[10]  | (\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )));
  assign new_n221_ = ~new_n220_ ^ (new_n176_ ^ ((~new_n179_ & (new_n117_ | (~new_n116_ & new_n125_) | (new_n116_ & ~new_n125_)) & (~new_n117_ | (~new_n116_ ^ new_n125_))) | (~new_n162_ & (new_n179_ | (~new_n117_ & (new_n116_ | ~new_n125_) & (~new_n116_ | new_n125_)) | (new_n117_ & (new_n116_ ^ new_n125_))) & (~new_n179_ | (~new_n117_ ^ (~new_n116_ ^ new_n125_))))));
  assign new_n222_ = (~new_n224_ | new_n242_) & ((~new_n225_ & (~new_n241_ | ((new_n244_ | (new_n223_ & ~new_n168_) | (~new_n223_ & new_n168_)) & (new_n227_ | (~new_n244_ & (~new_n223_ | new_n168_) & (new_n223_ | ~new_n168_)) | (new_n244_ & (~new_n223_ ^ ~new_n168_)))))) | (new_n224_ & ~new_n242_) | (~new_n224_ & new_n242_));
  assign new_n223_ = new_n167_ ^ ~new_n175_;
  assign new_n224_ = (new_n163_ ^ ~new_n164_) ^ ((new_n165_ & ~new_n166_) | (((~new_n167_ & new_n175_) | (~new_n168_ & (new_n167_ | ~new_n175_) & (~new_n167_ | new_n175_))) & (~new_n165_ | new_n166_) & (new_n165_ | ~new_n166_)));
  assign new_n225_ = ~new_n226_ & ((new_n165_ & ~new_n166_) | (~new_n165_ & new_n166_) | ((new_n167_ | ~new_n175_) & (new_n168_ | (~new_n167_ & new_n175_) | (new_n167_ & ~new_n175_)))) & ((new_n165_ ^ ~new_n166_) | (~new_n167_ & new_n175_) | (~new_n168_ & (new_n167_ | ~new_n175_) & (~new_n167_ | new_n175_)));
  assign new_n226_ = \a[29]  ^ ((((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))) | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & (~\b[8]  | (\a[26]  ^ \a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[9]  | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[7]  | (\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )));
  assign new_n227_ = (new_n228_ | ~new_n229_) & ((new_n228_ & ~new_n229_) | (~new_n228_ & new_n229_) | ((~new_n230_ | new_n231_) & (((new_n232_ | ~new_n240_) & (new_n233_ | (~new_n232_ & new_n240_) | (new_n232_ & ~new_n240_))) | (new_n230_ & ~new_n231_) | (~new_n230_ & new_n231_))));
  assign new_n228_ = \a[29]  ^ ((~new_n88_ | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & (~\b[6]  | (\a[26]  ^ \a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[7]  | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[5]  | (\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )));
  assign new_n229_ = (new_n172_ | (~new_n173_ & new_n174_)) ^ (new_n171_ ^ (~\a[32]  ^ (new_n170_ & (~new_n98_ | ~new_n169_))));
  assign new_n230_ = new_n173_ ^ ~new_n174_;
  assign new_n231_ = \a[29]  ^ ((~new_n91_ | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & (~\b[5]  | (\a[26]  ^ \a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[6]  | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[4]  | (\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )));
  assign new_n232_ = \a[29]  ^ ((~new_n94_ | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & (~\b[4]  | (\a[26]  ^ \a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[5]  | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[3]  | (\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )));
  assign new_n233_ = (~new_n236_ | (\a[29]  ^ (new_n235_ & (~new_n98_ | ~new_n234_)))) & ((~new_n237_ & (new_n238_ | ~new_n239_)) | (new_n236_ & (~\a[29]  ^ (new_n235_ & (~new_n98_ | ~new_n234_)))) | (~new_n236_ & (~\a[29]  | ~new_n235_ | (new_n98_ & new_n234_)) & (\a[29]  | (new_n235_ & (~new_n98_ | ~new_n234_)))));
  assign new_n234_ = (\a[26]  | \a[27] ) & (~\a[26]  | ~\a[27] ) & (~\a[28]  | ~\a[29] ) & (\a[28]  | \a[29] );
  assign new_n235_ = (~\b[3]  | (~\a[26]  ^ ~\a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[4]  | (~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[2]  | (\a[27]  ^ \a[28] ) | (~\a[26]  ^ ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] ));
  assign new_n236_ = ((\b[0]  & (\a[29]  ^ ~\a[30] ) & (~\a[30]  | ~\a[31] ) & (\a[30]  | \a[31] )) | (\b[1]  & (\a[29]  | \a[30] ) & (~\a[29]  | ~\a[30] ) & (~\a[31]  ^ \a[32] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & (\a[29]  | \a[30] ) & (~\a[29]  | ~\a[30] ) & (~\a[31]  | ~\a[32] ) & (\a[31]  | \a[32] ))) ^ (\a[32]  & \b[0]  & (\a[29]  | \a[30] ) & (~\a[29]  | ~\a[30] ));
  assign new_n237_ = \b[0]  & (~\a[29]  | ~\a[30] ) & (\a[29]  | \a[30] ) & (~\b[0]  | (~\a[26]  ^ ~\a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[1]  | (~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  ^ \a[29] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & \a[29]  & (~\b[0]  | (~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] )) & (~\b[0]  | (\a[27]  ^ \a[28] ) | (~\a[26]  ^ ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & (~\b[1]  | (~\a[26]  ^ ~\a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[2]  | (~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  ^ \a[29] )) & ((~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )));
  assign new_n238_ = \a[29]  ^ (((~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (~\a[26]  ^ ~\a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[3]  | (~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[1]  | (\a[27]  ^ \a[28] ) | (~\a[26]  ^ ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )));
  assign new_n239_ = (\b[0]  & (~\a[29]  | ~\a[30] ) & (\a[29]  | \a[30] )) ^ ((~\b[0]  | (~\a[26]  ^ ~\a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[1]  | (~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  ^ \a[29] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & \a[29]  & (~\b[0]  | (~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] )) & (~\b[0]  | (\a[27]  ^ \a[28] ) | (~\a[26]  ^ ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & (~\b[1]  | (~\a[26]  ^ ~\a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[2]  | (~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  ^ \a[29] )) & ((~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n240_ = (~\a[32]  | ((~\b[0]  | (~\a[29]  ^ ~\a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[1]  | (~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  ^ \a[32] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & \a[32]  & (~\b[0]  | (~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] )))) ^ ((~\b[1]  | (~\a[29]  ^ ~\a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[2]  | (~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  ^ \a[32] )) & ((~\a[29]  & ~\a[30] ) | (\a[29]  & \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (\a[30]  ^ \a[31] ) | (~\a[29]  ^ ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )));
  assign new_n241_ = ~new_n226_ ^ ((new_n165_ ^ ~new_n166_) ^ ((~new_n167_ & new_n175_) | (~new_n168_ & (new_n167_ | ~new_n175_) & (~new_n167_ | new_n175_))));
  assign new_n242_ = \a[29]  ^ (new_n243_ & (~new_n234_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n243_ = (~\b[9]  | (~\a[26]  ^ ~\a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[10]  | (~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[8]  | (\a[27]  ^ \a[28] ) | (~\a[26]  ^ ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] ));
  assign new_n244_ = \a[29]  ^ ((~\b[7]  | (\a[26]  ^ \a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[8]  | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[6]  | (\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & ((\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n79_ & (~\b[7]  ^ \b[8] ))));
  assign new_n245_ = ~new_n179_ ^ (~new_n117_ ^ (~new_n116_ ^ new_n125_));
  assign new_n246_ = \a[29]  ^ ((~new_n133_ | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & (~\b[12]  | (\a[26]  ^ \a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[13]  | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[11]  | (\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )));
  assign new_n247_ = \a[29]  ^ ((~new_n135_ | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & (~\b[10]  | (\a[26]  ^ \a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[11]  | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[9]  | (\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )));
  assign new_n248_ = new_n215_ & (~new_n180_ ^ (new_n211_ | (~new_n157_ & new_n212_)));
  assign new_n249_ = \a[29]  ^ ((~new_n186_ | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & (~\b[15]  | (\a[26]  ^ \a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[16]  | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[14]  | (\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )));
  assign new_n250_ = \a[29]  ^ ((~\b[13]  | (\a[26]  ^ \a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[14]  | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[12]  | (\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & ((\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n142_ & (~\b[13]  ^ \b[14] ))));
  assign new_n251_ = ~new_n208_ ^ (new_n184_ ^ (new_n204_ | (~new_n152_ & new_n205_)));
  assign new_n252_ = \a[29]  ^ ((~new_n253_ | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & (~\b[18]  | (\a[26]  ^ \a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[19]  | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[17]  | (\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )));
  assign new_n253_ = (\b[18]  ^ \b[19] ) ^ ((\b[17]  & \b[18] ) | ((~\b[17]  | ~\b[18] ) & (\b[17]  | \b[18] ) & ((\b[16]  & \b[17] ) | ((~\b[16]  | ~\b[17] ) & (\b[16]  | \b[17] ) & ((\b[15]  & \b[16] ) | ((~\b[15]  | ~\b[16] ) & (\b[15]  | \b[16] ) & ((\b[14]  & \b[15] ) | (((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] ))) & (~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] )))))))));
  assign new_n254_ = \a[29]  ^ ((~new_n144_ | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & (~\b[16]  | (\a[26]  ^ \a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[17]  | (\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  ^ \a[29] )) & (~\b[15]  | (\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )));
  assign new_n255_ = ~new_n200_ ^ (new_n189_ ^ (new_n74_ | (~new_n145_ & new_n188_)));
  assign new_n256_ = \a[29]  ^ (new_n258_ ^ (new_n257_ | (new_n189_ & (new_n74_ | (~new_n145_ & new_n188_)))));
  assign new_n257_ = ~new_n198_ & (~new_n191_ | (~new_n190_ & ~new_n197_)) & (new_n191_ | new_n190_ | new_n197_);
  assign new_n258_ = ~new_n265_ ^ (new_n260_ ^ (new_n259_ | (new_n191_ & (new_n190_ | new_n197_))));
  assign new_n259_ = ~new_n196_ & (~new_n192_ | new_n194_) & (new_n192_ | ~new_n194_);
  assign new_n260_ = ~new_n264_ ^ (new_n261_ ^ (new_n263_ | (new_n192_ & ~new_n194_)));
  assign new_n261_ = ~new_n262_ ^ (\a[38]  & ~\b[10] );
  assign new_n262_ = (~\b[11]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (\a[35]  ^ \a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[12]  | (\a[35]  ^ \a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[13]  | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  ^ \a[38] )) & (~new_n133_ | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ));
  assign new_n263_ = new_n193_ & \a[38]  & \b[9] ;
  assign new_n264_ = \a[35]  ^ ((~new_n186_ | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & (~\b[15]  | (\a[32]  ^ \a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[16]  | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[14]  | (\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )));
  assign new_n265_ = \a[32]  ^ ((~new_n253_ | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & (~\b[18]  | (\a[29]  ^ \a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[19]  | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  ^ \a[32] )) & (~\b[17]  | (\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )));
  assign new_n266_ = \a[29]  ^ (((\a[26]  & \a[27] ) | (~\a[26]  & ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] ) | (~new_n201_ ^ ~\b[19] )) & (~\b[19]  | (\a[26]  ^ \a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[18]  | (\a[27]  ^ \a[28] ) | (\a[26]  ^ \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )));
  assign new_n267_ = new_n255_ ^ ((~new_n266_ & (~new_n145_ | new_n188_) & (new_n145_ | ~new_n188_)) | (~new_n202_ & (new_n266_ | (new_n145_ & ~new_n188_) | (~new_n145_ & new_n188_)) & (~new_n266_ | (new_n145_ ^ ~new_n188_))));
  assign new_n268_ = (~new_n269_ | ~\a[26] ) & ((new_n269_ & \a[26] ) | (~new_n269_ & ~\a[26] ) | (~new_n273_ & (new_n273_ | new_n327_ | ((new_n328_ | (~new_n209_ & new_n271_) | (new_n209_ & ~new_n271_)) & (new_n275_ | (~new_n328_ & (new_n209_ | ~new_n271_) & (~new_n209_ | new_n271_)) | (new_n328_ & (new_n209_ ^ new_n271_)))))));
  assign new_n269_ = new_n272_ ^ (new_n207_ | (new_n251_ & (new_n270_ | (~new_n209_ & new_n271_))));
  assign new_n270_ = ~new_n254_ & (~new_n152_ | new_n205_) & (new_n152_ | ~new_n205_);
  assign new_n271_ = ~new_n254_ ^ (new_n152_ ^ ~new_n205_);
  assign new_n272_ = ~new_n252_ ^ (new_n206_ ^ (new_n150_ | (new_n184_ & (new_n204_ | (~new_n152_ & new_n205_)))));
  assign new_n273_ = ~new_n274_ & (~new_n251_ | (~new_n270_ & (new_n209_ | ~new_n271_))) & (new_n251_ | new_n270_ | (~new_n209_ & new_n271_));
  assign new_n274_ = \a[26]  ^ (~\b[19]  | (((\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & (new_n201_ | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ))));
  assign new_n275_ = (~new_n276_ | new_n324_) & ((new_n276_ & ~new_n324_) | (~new_n276_ & new_n324_) | ((~new_n278_ | new_n325_) & ((new_n278_ & ~new_n325_) | (~new_n278_ & new_n325_) | ((new_n326_ | (~new_n216_ & new_n323_) | (new_n216_ & ~new_n323_)) & (new_n279_ | (~new_n326_ & (new_n216_ | ~new_n323_) & (~new_n216_ | new_n323_)) | (new_n326_ & (new_n216_ ^ new_n323_)))))));
  assign new_n276_ = new_n277_ ^ (new_n214_ | (((~new_n250_ & (new_n157_ | ~new_n212_) & (~new_n157_ | new_n212_)) | (~new_n216_ & (new_n250_ | (~new_n157_ & new_n212_) | (new_n157_ & ~new_n212_)) & (~new_n250_ | (~new_n157_ ^ new_n212_)))) & ~new_n214_ & ~new_n248_));
  assign new_n277_ = ~new_n249_ ^ (new_n213_ ^ (new_n155_ | (new_n180_ & (new_n211_ | (~new_n157_ & new_n212_)))));
  assign new_n278_ = (~new_n214_ & ~new_n248_) ^ ((~new_n250_ & (new_n157_ | ~new_n212_) & (~new_n157_ | new_n212_)) | (~new_n216_ & (new_n250_ | (~new_n157_ & new_n212_) | (new_n157_ & ~new_n212_)) & (~new_n250_ | (~new_n157_ ^ new_n212_))));
  assign new_n279_ = (~new_n280_ | new_n321_) & ((new_n280_ & ~new_n321_) | (~new_n280_ & new_n321_) | (~new_n284_ & (new_n284_ | new_n320_ | ((new_n322_ | (~new_n222_ & new_n282_) | (new_n222_ & ~new_n282_)) & (new_n286_ | (~new_n322_ & (new_n222_ | ~new_n282_) & (~new_n222_ | new_n282_)) | (new_n322_ & (new_n222_ ^ new_n282_)))))));
  assign new_n280_ = new_n283_ ^ (new_n219_ | (new_n221_ & (new_n281_ | (~new_n222_ & new_n282_))));
  assign new_n281_ = ~new_n247_ & (~new_n162_ | new_n245_) & (new_n162_ | ~new_n245_);
  assign new_n282_ = ~new_n247_ ^ (new_n162_ ^ ~new_n245_);
  assign new_n283_ = ~new_n246_ ^ (new_n218_ ^ (new_n160_ | (new_n176_ & ((~new_n179_ & (~new_n158_ | new_n117_) & (new_n158_ | ~new_n117_)) | (~new_n162_ & (new_n179_ | (new_n158_ & ~new_n117_) | (~new_n158_ & new_n117_)) & (~new_n179_ | (new_n158_ ^ ~new_n117_)))))));
  assign new_n284_ = ~new_n285_ & (~new_n221_ | (~new_n281_ & (new_n222_ | ~new_n282_))) & (new_n221_ | new_n281_ | (~new_n222_ & new_n282_));
  assign new_n285_ = \a[26]  ^ ((((~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] ) & ((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )))) | ((~\b[14]  ^ \b[15] ) & (~\b[13]  | ~\b[14] ) & (new_n142_ | (\b[13]  & \b[14] ) | (~\b[13]  & ~\b[14] ))) | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & (~\b[14]  | (\a[23]  ^ \a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[15]  | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[13]  | (\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )));
  assign new_n286_ = (~new_n287_ | new_n319_) & ((new_n287_ & ~new_n319_) | (~new_n287_ & new_n319_) | (~new_n289_ & (~new_n291_ | (~new_n292_ & (new_n295_ | ~new_n318_)))));
  assign new_n287_ = new_n288_ ^ (new_n225_ | (new_n241_ & ((~new_n244_ & (new_n168_ | (~new_n167_ & new_n175_) | (new_n167_ & ~new_n175_)) & (~new_n168_ | (~new_n167_ ^ new_n175_))) | (~new_n227_ & (new_n244_ | (~new_n168_ & (new_n167_ | ~new_n175_) & (~new_n167_ | new_n175_)) | (new_n168_ & (new_n167_ ^ new_n175_))) & (~new_n244_ | (~new_n168_ ^ (~new_n167_ ^ new_n175_)))))));
  assign new_n288_ = ~new_n242_ ^ ((new_n163_ ^ ~new_n164_) ^ ((new_n165_ & ~new_n166_) | ((~new_n165_ | new_n166_) & (new_n165_ | ~new_n166_) & ((~new_n167_ & new_n175_) | (~new_n168_ & (new_n167_ | ~new_n175_) & (~new_n167_ | new_n175_))))));
  assign new_n289_ = ~new_n290_ & (~new_n241_ | ((new_n244_ | (~new_n168_ & (new_n167_ | ~new_n175_) & (~new_n167_ | new_n175_)) | (new_n168_ & (new_n167_ ^ new_n175_))) & (new_n227_ | (~new_n244_ & (new_n168_ | (~new_n167_ & new_n175_) | (new_n167_ & ~new_n175_)) & (~new_n168_ | (~new_n167_ ^ new_n175_))) | (new_n244_ & (new_n168_ ^ (~new_n167_ ^ new_n175_)))))) & (new_n241_ | (~new_n244_ & (new_n168_ | (~new_n167_ & new_n175_) | (new_n167_ & ~new_n175_)) & (~new_n168_ | (~new_n167_ ^ new_n175_))) | (~new_n227_ & (new_n244_ | (~new_n168_ & (new_n167_ | ~new_n175_) & (~new_n167_ | new_n175_)) | (new_n168_ & (new_n167_ ^ new_n175_))) & (~new_n244_ | (~new_n168_ ^ (~new_n167_ ^ new_n175_)))));
  assign new_n290_ = \a[26]  ^ ((~new_n107_ | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & (~\b[11]  | (\a[23]  ^ \a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[12]  | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[10]  | (\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )));
  assign new_n291_ = ~new_n290_ ^ (new_n241_ ^ ((~new_n244_ & (new_n168_ | (~new_n167_ & new_n175_) | (new_n167_ & ~new_n175_)) & (~new_n168_ | (~new_n167_ ^ new_n175_))) | (~new_n227_ & (new_n244_ | (~new_n168_ & (new_n167_ | ~new_n175_) & (~new_n167_ | new_n175_)) | (new_n168_ & (new_n167_ ^ new_n175_))) & (~new_n244_ | (~new_n168_ ^ (~new_n167_ ^ new_n175_))))));
  assign new_n292_ = ~new_n294_ & (~new_n227_ | new_n293_) & (new_n227_ | ~new_n293_);
  assign new_n293_ = ~new_n244_ ^ (~new_n168_ ^ (~new_n167_ ^ new_n175_));
  assign new_n294_ = \a[26]  ^ ((~new_n135_ | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & (~\b[10]  | (\a[23]  ^ \a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[11]  | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[9]  | (\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )));
  assign new_n295_ = (~new_n297_ | new_n315_) & ((~new_n298_ & (~new_n314_ | ((new_n317_ | (new_n296_ & ~new_n233_) | (~new_n296_ & new_n233_)) & (new_n300_ | (~new_n317_ & (~new_n296_ | new_n233_) & (new_n296_ | ~new_n233_)) | (new_n317_ & (~new_n296_ ^ ~new_n233_)))))) | (new_n297_ & ~new_n315_) | (~new_n297_ & new_n315_));
  assign new_n296_ = new_n232_ ^ ~new_n240_;
  assign new_n297_ = (new_n228_ ^ ~new_n229_) ^ ((new_n230_ & ~new_n231_) | (((~new_n232_ & new_n240_) | (~new_n233_ & (new_n232_ | ~new_n240_) & (~new_n232_ | new_n240_))) & (~new_n230_ | new_n231_) & (new_n230_ | ~new_n231_)));
  assign new_n298_ = ~new_n299_ & ((new_n230_ & ~new_n231_) | (~new_n230_ & new_n231_) | ((new_n232_ | ~new_n240_) & (new_n233_ | (~new_n232_ & new_n240_) | (new_n232_ & ~new_n240_)))) & ((new_n230_ ^ ~new_n231_) | (~new_n232_ & new_n240_) | (~new_n233_ & (new_n232_ | ~new_n240_) & (~new_n232_ | new_n240_)));
  assign new_n299_ = \a[26]  ^ ((((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))) | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & (~\b[8]  | (\a[23]  ^ \a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[9]  | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[7]  | (\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )));
  assign new_n300_ = (new_n301_ | ~new_n302_) & ((new_n301_ & ~new_n302_) | (~new_n301_ & new_n302_) | ((~new_n303_ | new_n304_) & (((new_n305_ | ~new_n313_) & (new_n306_ | (~new_n305_ & new_n313_) | (new_n305_ & ~new_n313_))) | (new_n303_ & ~new_n304_) | (~new_n303_ & new_n304_))));
  assign new_n301_ = \a[26]  ^ ((~new_n88_ | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & (~\b[6]  | (\a[23]  ^ \a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[7]  | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[5]  | (\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )));
  assign new_n302_ = (new_n237_ | (~new_n238_ & new_n239_)) ^ (new_n236_ ^ (~\a[29]  ^ (new_n235_ & (~new_n98_ | ~new_n234_))));
  assign new_n303_ = new_n238_ ^ ~new_n239_;
  assign new_n304_ = \a[26]  ^ ((~new_n91_ | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & (~\b[5]  | (\a[23]  ^ \a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[6]  | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[4]  | (\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )));
  assign new_n305_ = \a[26]  ^ ((~new_n94_ | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & (~\b[4]  | (\a[23]  ^ \a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[5]  | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[3]  | (\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )));
  assign new_n306_ = (~new_n309_ | (\a[26]  ^ (new_n308_ & (~new_n98_ | ~new_n307_)))) & ((~new_n310_ & (new_n311_ | ~new_n312_)) | (new_n309_ & (~\a[26]  ^ (new_n308_ & (~new_n98_ | ~new_n307_)))) | (~new_n309_ & (~\a[26]  | ~new_n308_ | (new_n98_ & new_n307_)) & (\a[26]  | (new_n308_ & (~new_n98_ | ~new_n307_)))));
  assign new_n307_ = (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] ) & (~\a[25]  | ~\a[26] ) & (\a[25]  | \a[26] );
  assign new_n308_ = (~\b[3]  | (~\a[23]  ^ ~\a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[4]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[2]  | (\a[24]  ^ \a[25] ) | (~\a[23]  ^ ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ));
  assign new_n309_ = ((\b[0]  & (\a[26]  ^ ~\a[27] ) & (~\a[27]  | ~\a[28] ) & (\a[27]  | \a[28] )) | (\b[1]  & (\a[26]  | \a[27] ) & (~\a[26]  | ~\a[27] ) & (~\a[28]  ^ \a[29] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & (\a[26]  | \a[27] ) & (~\a[26]  | ~\a[27] ) & (~\a[28]  | ~\a[29] ) & (\a[28]  | \a[29] ))) ^ (\a[29]  & \b[0]  & (\a[26]  | \a[27] ) & (~\a[26]  | ~\a[27] ));
  assign new_n310_ = \b[0]  & (~\a[26]  | ~\a[27] ) & (\a[26]  | \a[27] ) & (~\b[0]  | (~\a[23]  ^ ~\a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[1]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  ^ \a[26] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & \a[26]  & (~\b[0]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~\b[0]  | (\a[24]  ^ \a[25] ) | (~\a[23]  ^ ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & (~\b[1]  | (~\a[23]  ^ ~\a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[2]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  ^ \a[26] )) & ((~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )));
  assign new_n311_ = \a[26]  ^ (((~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (~\a[23]  ^ ~\a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[3]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[1]  | (\a[24]  ^ \a[25] ) | (~\a[23]  ^ ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )));
  assign new_n312_ = (\b[0]  & (~\a[26]  | ~\a[27] ) & (\a[26]  | \a[27] )) ^ ((~\b[0]  | (~\a[23]  ^ ~\a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[1]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  ^ \a[26] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & \a[26]  & (~\b[0]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )) & (~\b[0]  | (\a[24]  ^ \a[25] ) | (~\a[23]  ^ ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & (~\b[1]  | (~\a[23]  ^ ~\a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[2]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  ^ \a[26] )) & ((~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n313_ = (~\a[29]  | ((~\b[0]  | (~\a[26]  ^ ~\a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[1]  | (~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  ^ \a[29] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )) & \a[29]  & (~\b[0]  | (~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] )))) ^ ((~\b[1]  | (~\a[26]  ^ ~\a[27] ) | (\a[27]  & \a[28] ) | (~\a[27]  & ~\a[28] )) & (~\b[2]  | (~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  ^ \a[29] )) & ((~\a[26]  & ~\a[27] ) | (\a[26]  & \a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (\a[27]  ^ \a[28] ) | (~\a[26]  ^ ~\a[27] ) | (\a[28]  & \a[29] ) | (~\a[28]  & ~\a[29] )));
  assign new_n314_ = ~new_n299_ ^ ((new_n230_ ^ ~new_n231_) ^ ((~new_n232_ & new_n240_) | (~new_n233_ & (new_n232_ | ~new_n240_) & (~new_n232_ | new_n240_))));
  assign new_n315_ = \a[26]  ^ (new_n316_ & (~new_n307_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n316_ = (~\b[9]  | (~\a[23]  ^ ~\a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[10]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[8]  | (\a[24]  ^ \a[25] ) | (~\a[23]  ^ ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ));
  assign new_n317_ = \a[26]  ^ ((~\b[7]  | (\a[23]  ^ \a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[8]  | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[6]  | (\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & ((\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n79_ & (~\b[7]  ^ \b[8] ))));
  assign new_n318_ = ~new_n294_ ^ (new_n227_ ^ ~new_n293_);
  assign new_n319_ = \a[26]  ^ ((~new_n133_ | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & (~\b[12]  | (\a[23]  ^ \a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[13]  | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[11]  | (\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )));
  assign new_n320_ = new_n285_ & (~new_n221_ ^ (new_n281_ | (~new_n222_ & new_n282_)));
  assign new_n321_ = \a[26]  ^ ((~new_n186_ | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & (~\b[15]  | (\a[23]  ^ \a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[16]  | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[14]  | (\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )));
  assign new_n322_ = \a[26]  ^ ((~\b[13]  | (\a[23]  ^ \a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[14]  | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[12]  | (\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & ((\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n142_ & (~\b[13]  ^ \b[14] ))));
  assign new_n323_ = ~new_n250_ ^ (new_n157_ ^ ~new_n212_);
  assign new_n324_ = \a[26]  ^ ((~new_n253_ | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & (~\b[18]  | (\a[23]  ^ \a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[19]  | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[17]  | (\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )));
  assign new_n325_ = \a[26]  ^ ((~new_n199_ | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & (~\b[17]  | (\a[23]  ^ \a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[18]  | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[16]  | (\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )));
  assign new_n326_ = \a[26]  ^ ((~new_n144_ | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & (~\b[16]  | (\a[23]  ^ \a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[17]  | (\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  ^ \a[26] )) & (~\b[15]  | (\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )));
  assign new_n327_ = new_n274_ & (~new_n251_ ^ (new_n270_ | (~new_n209_ & new_n271_)));
  assign new_n328_ = \a[26]  ^ (((\a[23]  & \a[24] ) | (~\a[23]  & ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (~new_n201_ ^ ~\b[19] )) & (~\b[19]  | (\a[23]  ^ \a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[18]  | (\a[24]  ^ \a[25] ) | (\a[23]  ^ \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )));
  assign new_n329_ = ~new_n266_ ^ (new_n145_ ^ ~new_n188_);
  assign new_n330_ = \a[26]  ^ (new_n331_ ^ ~new_n333_);
  assign new_n331_ = (~new_n332_ | ~\a[29] ) & ((new_n332_ & \a[29] ) | (~new_n332_ & ~\a[29] ) | (~new_n73_ & (~new_n255_ | ((new_n266_ | (~new_n145_ & new_n188_) | (new_n145_ & ~new_n188_)) & (new_n202_ | (~new_n266_ & (new_n145_ | ~new_n188_) & (~new_n145_ | new_n188_)) | (new_n266_ & (new_n145_ ^ new_n188_)))))));
  assign new_n332_ = new_n258_ ^ (new_n257_ | (new_n189_ & (new_n74_ | (~new_n145_ & new_n188_))));
  assign new_n333_ = ~new_n334_ ^ ~\a[29] ;
  assign new_n334_ = new_n336_ ^ ((new_n335_ & ~new_n265_) | ((new_n257_ | (new_n189_ & (new_n74_ | (~new_n145_ & new_n188_)))) & (~new_n335_ | new_n265_) & (new_n335_ | ~new_n265_)));
  assign new_n335_ = new_n260_ ^ (new_n259_ | (new_n191_ & (new_n190_ | new_n197_)));
  assign new_n336_ = ~new_n343_ ^ (new_n338_ ^ (new_n337_ | (new_n260_ & (new_n259_ | (new_n191_ & (new_n190_ | new_n197_))))));
  assign new_n337_ = ~new_n264_ & (~new_n261_ | (~new_n263_ & (~new_n192_ | new_n194_))) & (new_n261_ | new_n263_ | (new_n192_ & ~new_n194_));
  assign new_n338_ = ~new_n339_ ^ (new_n340_ ^ (new_n342_ | (new_n261_ & (new_n263_ | (new_n192_ & ~new_n194_)))));
  assign new_n339_ = \a[35]  ^ ((~new_n144_ | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & (~\b[16]  | (\a[32]  ^ \a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[17]  | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[15]  | (\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )));
  assign new_n340_ = ~new_n341_ ^ (\a[38]  & ~\b[11] );
  assign new_n341_ = (~\b[12]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (\a[35]  ^ \a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[13]  | (\a[35]  ^ \a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[14]  | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  ^ \a[38] )) & ((\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n142_ & (~\b[13]  ^ \b[14] )));
  assign new_n342_ = new_n262_ & \a[38]  & \b[10] ;
  assign new_n343_ = \a[32]  ^ (((\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] ) | (~new_n201_ ^ ~\b[19] )) & (~\b[19]  | (\a[29]  ^ \a[30] ) | (\a[30]  & \a[31] ) | (~\a[30]  & ~\a[31] )) & (~\b[18]  | (\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )));
  assign new_n344_ = ((\a[23]  & (~new_n71_ | new_n330_) & (new_n71_ | ~new_n330_)) | ((~\a[23]  | (new_n71_ & ~new_n330_) | (~new_n71_ & new_n330_)) & (\a[23]  | (new_n71_ ^ ~new_n330_)) & ((new_n361_ & \a[23] ) | ((~new_n361_ | ~\a[23] ) & (new_n361_ | \a[23] ) & ((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] ))))))) ^ (\a[23]  ^ (new_n345_ ^ ~new_n346_));
  assign new_n345_ = (~\a[26]  | (new_n331_ & ~new_n333_) | (~new_n331_ & new_n333_)) & ((\a[26]  & (~new_n331_ | new_n333_) & (new_n331_ | ~new_n333_)) | (~\a[26]  & (~new_n331_ ^ ~new_n333_)) | ((~new_n72_ | ~\a[26] ) & ((new_n72_ & \a[26] ) | (~new_n72_ & ~\a[26] ) | ((~new_n267_ | ~\a[26] ) & ((new_n267_ & \a[26] ) | (~new_n267_ & ~\a[26] ) | ((~\a[26]  | (~new_n202_ & new_n329_) | (new_n202_ & ~new_n329_)) & (new_n268_ | (\a[26]  & (new_n202_ | ~new_n329_) & (~new_n202_ | new_n329_)) | (~\a[26]  & (new_n202_ ^ new_n329_)))))))));
  assign new_n346_ = \a[26]  ^ (((new_n334_ & \a[29] ) | (~new_n331_ & (~new_n334_ | ~\a[29] ) & (new_n334_ | \a[29] ))) ^ (~new_n347_ ^ ~\a[29] ));
  assign new_n347_ = new_n349_ ^ (new_n348_ | new_n360_);
  assign new_n348_ = new_n336_ & ((new_n335_ & ~new_n265_) | ((new_n257_ | (new_n189_ & (new_n74_ | (~new_n145_ & new_n188_)))) & (~new_n335_ | new_n265_) & (new_n335_ | ~new_n265_)));
  assign new_n349_ = ~new_n359_ ^ (new_n350_ ^ ~new_n352_);
  assign new_n350_ = (~new_n351_ | new_n339_) & ((~new_n337_ & (~new_n260_ | (~new_n259_ & (~new_n191_ | (~new_n190_ & ~new_n197_))))) | (new_n351_ & ~new_n339_) | (~new_n351_ & new_n339_));
  assign new_n351_ = new_n340_ ^ (new_n342_ | (new_n261_ & (new_n263_ | (new_n192_ & ~new_n194_))));
  assign new_n352_ = ~new_n354_ ^ (new_n355_ ^ (new_n358_ | (~new_n353_ & new_n340_)));
  assign new_n353_ = ~new_n342_ & (~new_n261_ | (~new_n263_ & (~new_n192_ | new_n194_)));
  assign new_n354_ = \a[35]  ^ ((~new_n199_ | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & (~\b[17]  | (\a[32]  ^ \a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[18]  | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[16]  | (\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )));
  assign new_n355_ = (\a[38]  & ~\b[12] ) ^ (~new_n357_ | (new_n356_ & new_n80_));
  assign new_n356_ = ((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] ))) ^ (\b[14]  ^ \b[15] );
  assign new_n357_ = (~\b[13]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (~\a[35]  ^ ~\a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[14]  | (~\a[35]  ^ ~\a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[15]  | (~\a[35]  & ~\a[36] ) | (\a[35]  & \a[36] ) | (\a[37]  ^ \a[38] ));
  assign new_n358_ = new_n341_ & \a[38]  & \b[11] ;
  assign new_n359_ = \a[32]  ^ (~\b[19]  | (((\a[30]  ^ \a[31] ) | (\a[29]  ^ \a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] )) & (new_n201_ | (\a[29]  & \a[30] ) | (~\a[29]  & ~\a[30] ) | (\a[31]  & \a[32] ) | (~\a[31]  & ~\a[32] ))));
  assign new_n360_ = ~new_n343_ & (~new_n338_ | (~new_n337_ & (~new_n260_ | (~new_n259_ & (~new_n191_ | (~new_n190_ & ~new_n197_)))))) & (new_n338_ | new_n337_ | (new_n260_ & (new_n259_ | (new_n191_ & (new_n190_ | new_n197_)))));
  assign new_n361_ = ((new_n267_ & \a[26] ) | ((~new_n267_ | ~\a[26] ) & (new_n267_ | \a[26] ) & ((\a[26]  & (new_n202_ | ~new_n329_) & (~new_n202_ | new_n329_)) | (~new_n268_ & (~\a[26]  | (~new_n202_ & new_n329_) | (new_n202_ & ~new_n329_)) & (\a[26]  | (~new_n202_ ^ new_n329_)))))) ^ (new_n72_ ^ \a[26] );
  assign new_n362_ = ((\a[26]  & (~new_n202_ | new_n329_) & (new_n202_ | ~new_n329_)) | (~new_n268_ & (~\a[26]  | (new_n202_ & ~new_n329_) | (~new_n202_ & new_n329_)) & (\a[26]  | (new_n202_ ^ ~new_n329_)))) ^ (new_n267_ ^ \a[26] );
  assign new_n363_ = (~\a[23]  | (new_n268_ & ~new_n364_) | (~new_n268_ & new_n364_)) & (((~new_n365_ | ~\a[23] ) & ((new_n365_ & \a[23] ) | (~new_n365_ & ~\a[23] ) | ((~new_n367_ | ~\a[23] ) & (((~new_n368_ | ~\a[23] ) & (new_n370_ | (~new_n368_ & ~\a[23] ) | (new_n368_ & \a[23] ))) | (new_n367_ & \a[23] ) | (~new_n367_ & ~\a[23] ))))) | (\a[23]  & (~new_n268_ | new_n364_) & (new_n268_ | ~new_n364_)) | (~\a[23]  & (~new_n268_ ^ ~new_n364_)));
  assign new_n364_ = \a[26]  ^ (new_n202_ ^ ~new_n329_);
  assign new_n365_ = new_n366_ ^ (new_n273_ | (((~new_n328_ & (new_n209_ | ~new_n271_) & (~new_n209_ | new_n271_)) | (~new_n275_ & (new_n328_ | (~new_n209_ & new_n271_) | (new_n209_ & ~new_n271_)) & (~new_n328_ | (~new_n209_ ^ new_n271_)))) & ~new_n273_ & ~new_n327_));
  assign new_n366_ = \a[26]  ^ (new_n272_ ^ (new_n207_ | (new_n251_ & (new_n270_ | (~new_n209_ & new_n271_)))));
  assign new_n367_ = (~new_n273_ & ~new_n327_) ^ ((~new_n328_ & (new_n209_ | ~new_n271_) & (~new_n209_ | new_n271_)) | (~new_n275_ & (new_n328_ | (~new_n209_ & new_n271_) | (new_n209_ & ~new_n271_)) & (~new_n328_ | (~new_n209_ ^ new_n271_))));
  assign new_n368_ = new_n275_ ^ ~new_n369_;
  assign new_n369_ = ~new_n328_ ^ (new_n209_ ^ ~new_n271_);
  assign new_n370_ = (~new_n371_ | ~\a[23] ) & ((new_n371_ & \a[23] ) | (~new_n371_ & ~\a[23] ) | (~new_n372_ & (~new_n426_ | ((new_n428_ | (~new_n279_ & new_n427_) | (new_n279_ & ~new_n427_)) & (new_n374_ | (~new_n428_ & (new_n279_ | ~new_n427_) & (~new_n279_ | new_n427_)) | (new_n428_ & (new_n279_ ^ new_n427_)))))));
  assign new_n371_ = (new_n276_ ^ ~new_n324_) ^ ((new_n278_ & ~new_n325_) | ((~new_n278_ | new_n325_) & (new_n278_ | ~new_n325_) & ((~new_n326_ & (new_n216_ | ~new_n323_) & (~new_n216_ | new_n323_)) | (~new_n279_ & (new_n326_ | (~new_n216_ & new_n323_) | (new_n216_ & ~new_n323_)) & (~new_n326_ | (~new_n216_ ^ new_n323_))))));
  assign new_n372_ = ~new_n373_ & ((~new_n278_ & new_n325_) | (new_n278_ & ~new_n325_) | ((new_n326_ | (new_n216_ & ~new_n323_) | (~new_n216_ & new_n323_)) & (new_n279_ | (~new_n326_ & (~new_n216_ | new_n323_) & (new_n216_ | ~new_n323_)) | (new_n326_ & (~new_n216_ ^ ~new_n323_))))) & ((~new_n278_ ^ new_n325_) | (~new_n326_ & (~new_n216_ | new_n323_) & (new_n216_ | ~new_n323_)) | (~new_n279_ & (new_n326_ | (new_n216_ & ~new_n323_) | (~new_n216_ & new_n323_)) & (~new_n326_ | (new_n216_ ^ ~new_n323_))));
  assign new_n373_ = \a[23]  ^ (~\b[19]  | (((\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (new_n201_ | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ))));
  assign new_n374_ = (~new_n375_ | new_n425_) & ((new_n375_ & ~new_n425_) | (~new_n375_ & new_n425_) | (~new_n377_ & (~new_n424_ | (~new_n379_ & (new_n382_ | ~new_n423_)))));
  assign new_n375_ = new_n376_ ^ (new_n284_ | (((~new_n322_ & (new_n222_ | ~new_n282_) & (~new_n222_ | new_n282_)) | (~new_n286_ & (new_n322_ | (~new_n222_ & new_n282_) | (new_n222_ & ~new_n282_)) & (~new_n322_ | (~new_n222_ ^ new_n282_)))) & ~new_n284_ & ~new_n320_));
  assign new_n376_ = ~new_n321_ ^ (new_n283_ ^ (new_n219_ | (new_n221_ & (new_n281_ | (~new_n222_ & new_n282_)))));
  assign new_n377_ = ~new_n378_ & (new_n284_ | new_n320_ | ((new_n322_ | (~new_n222_ & new_n282_) | (new_n222_ & ~new_n282_)) & (new_n286_ | (~new_n322_ & (new_n222_ | ~new_n282_) & (~new_n222_ | new_n282_)) | (new_n322_ & (new_n222_ ^ new_n282_))))) & ((~new_n284_ & ~new_n320_) | (~new_n322_ & (new_n222_ | ~new_n282_) & (~new_n222_ | new_n282_)) | (~new_n286_ & (new_n322_ | (~new_n222_ & new_n282_) | (new_n222_ & ~new_n282_)) & (~new_n322_ | (~new_n222_ ^ new_n282_))));
  assign new_n378_ = \a[23]  ^ ((~\b[16]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[17]  | (\a[20]  ^ \a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[18]  | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  ^ \a[23] )) & (~new_n199_ | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] )));
  assign new_n379_ = ~new_n381_ & (~new_n286_ | new_n380_) & (new_n286_ | ~new_n380_);
  assign new_n380_ = ~new_n322_ ^ (new_n222_ ^ ~new_n282_);
  assign new_n381_ = \a[23]  ^ ((~\b[15]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[16]  | (\a[20]  ^ \a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[17]  | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  ^ \a[23] )) & (~new_n144_ | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] )));
  assign new_n382_ = (~new_n383_ | new_n421_) & ((new_n383_ & ~new_n421_) | (~new_n383_ & new_n421_) | (~new_n384_ & (new_n384_ | new_n420_ | ((new_n422_ | (~new_n295_ & new_n318_) | (new_n295_ & ~new_n318_)) & (new_n386_ | (~new_n422_ & (new_n295_ | ~new_n318_) & (~new_n295_ | new_n318_)) | (new_n422_ & (new_n295_ ^ new_n318_)))))));
  assign new_n383_ = (new_n287_ ^ ~new_n319_) ^ (new_n289_ | (new_n291_ & (new_n292_ | (~new_n295_ & new_n318_))));
  assign new_n384_ = ~new_n385_ & (~new_n291_ | (~new_n292_ & (new_n295_ | ~new_n318_))) & (new_n291_ | new_n292_ | (~new_n295_ & new_n318_));
  assign new_n385_ = \a[23]  ^ ((((~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] ) & ((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )))) | ((~\b[14]  ^ \b[15] ) & (~\b[13]  | ~\b[14] ) & (new_n142_ | (\b[13]  & \b[14] ) | (~\b[13]  & ~\b[14] ))) | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] )) & (~\b[13]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[14]  | (\a[20]  ^ \a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[15]  | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  ^ \a[23] )));
  assign new_n386_ = (~new_n387_ | new_n419_) & ((new_n387_ & ~new_n419_) | (~new_n387_ & new_n419_) | (~new_n389_ & (~new_n418_ | (~new_n391_ & (new_n394_ | ~new_n417_)))));
  assign new_n387_ = new_n388_ ^ (new_n298_ | (new_n314_ & ((~new_n317_ & (new_n233_ | (~new_n232_ & new_n240_) | (new_n232_ & ~new_n240_)) & (~new_n233_ | (~new_n232_ ^ new_n240_))) | (~new_n300_ & (new_n317_ | (~new_n233_ & (new_n232_ | ~new_n240_) & (~new_n232_ | new_n240_)) | (new_n233_ & (new_n232_ ^ new_n240_))) & (~new_n317_ | (~new_n233_ ^ (~new_n232_ ^ new_n240_)))))));
  assign new_n388_ = ~new_n315_ ^ ((new_n228_ ^ ~new_n229_) ^ ((new_n230_ & ~new_n231_) | ((~new_n230_ | new_n231_) & (new_n230_ | ~new_n231_) & ((~new_n232_ & new_n240_) | (~new_n233_ & (new_n232_ | ~new_n240_) & (~new_n232_ | new_n240_))))));
  assign new_n389_ = ~new_n390_ & (~new_n314_ | ((new_n317_ | (~new_n233_ & (new_n232_ | ~new_n240_) & (~new_n232_ | new_n240_)) | (new_n233_ & (new_n232_ ^ new_n240_))) & (new_n300_ | (~new_n317_ & (new_n233_ | (~new_n232_ & new_n240_) | (new_n232_ & ~new_n240_)) & (~new_n233_ | (~new_n232_ ^ new_n240_))) | (new_n317_ & (new_n233_ ^ (~new_n232_ ^ new_n240_)))))) & (new_n314_ | (~new_n317_ & (new_n233_ | (~new_n232_ & new_n240_) | (new_n232_ & ~new_n240_)) & (~new_n233_ | (~new_n232_ ^ new_n240_))) | (~new_n300_ & (new_n317_ | (~new_n233_ & (new_n232_ | ~new_n240_) & (~new_n232_ | new_n240_)) | (new_n233_ & (new_n232_ ^ new_n240_))) & (~new_n317_ | (~new_n233_ ^ (~new_n232_ ^ new_n240_)))));
  assign new_n390_ = \a[23]  ^ ((~\b[10]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[11]  | (\a[20]  ^ \a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[12]  | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  ^ \a[23] )) & (~new_n107_ | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] )));
  assign new_n391_ = ~new_n393_ & (~new_n300_ | new_n392_) & (new_n300_ | ~new_n392_);
  assign new_n392_ = ~new_n317_ ^ (~new_n233_ ^ (~new_n232_ ^ new_n240_));
  assign new_n393_ = \a[23]  ^ ((~\b[9]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[10]  | (\a[20]  ^ \a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[11]  | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  ^ \a[23] )) & (~new_n135_ | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] )));
  assign new_n394_ = (~new_n396_ | new_n414_) & ((~new_n397_ & (~new_n413_ | ((new_n416_ | (new_n395_ & ~new_n306_) | (~new_n395_ & new_n306_)) & (new_n399_ | (~new_n416_ & (~new_n395_ | new_n306_) & (new_n395_ | ~new_n306_)) | (new_n416_ & (~new_n395_ ^ ~new_n306_)))))) | (new_n396_ & ~new_n414_) | (~new_n396_ & new_n414_));
  assign new_n395_ = new_n305_ ^ ~new_n313_;
  assign new_n396_ = (new_n301_ ^ ~new_n302_) ^ ((new_n303_ & ~new_n304_) | (((~new_n305_ & new_n313_) | (~new_n306_ & (new_n305_ | ~new_n313_) & (~new_n305_ | new_n313_))) & (~new_n303_ | new_n304_) & (new_n303_ | ~new_n304_)));
  assign new_n397_ = ~new_n398_ & ((new_n303_ & ~new_n304_) | (~new_n303_ & new_n304_) | ((new_n305_ | ~new_n313_) & (new_n306_ | (~new_n305_ & new_n313_) | (new_n305_ & ~new_n313_)))) & ((new_n303_ ^ ~new_n304_) | (~new_n305_ & new_n313_) | (~new_n306_ & (new_n305_ | ~new_n313_) & (~new_n305_ | new_n313_)));
  assign new_n398_ = \a[23]  ^ ((((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))) | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] )) & (~\b[7]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[8]  | (\a[20]  ^ \a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[9]  | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  ^ \a[23] )));
  assign new_n399_ = (new_n400_ | ~new_n401_) & ((new_n400_ & ~new_n401_) | (~new_n400_ & new_n401_) | ((~new_n402_ | new_n403_) & (((new_n404_ | ~new_n412_) & (new_n405_ | (~new_n404_ & new_n412_) | (new_n404_ & ~new_n412_))) | (new_n402_ & ~new_n403_) | (~new_n402_ & new_n403_))));
  assign new_n400_ = \a[23]  ^ ((~\b[5]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[6]  | (\a[20]  ^ \a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[7]  | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  ^ \a[23] )) & (~new_n88_ | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] )));
  assign new_n401_ = (new_n310_ | (~new_n311_ & new_n312_)) ^ (new_n309_ ^ (~\a[26]  ^ (new_n308_ & (~new_n98_ | ~new_n307_))));
  assign new_n402_ = new_n311_ ^ ~new_n312_;
  assign new_n403_ = \a[23]  ^ ((~\b[4]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[5]  | (\a[20]  ^ \a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[6]  | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  ^ \a[23] )) & (~new_n91_ | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] )));
  assign new_n404_ = \a[23]  ^ ((~\b[3]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[4]  | (\a[20]  ^ \a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[5]  | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  ^ \a[23] )) & (~new_n94_ | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] )));
  assign new_n405_ = (~new_n408_ | (\a[23]  ^ (new_n407_ & (~new_n98_ | ~new_n406_)))) & ((~new_n409_ & (new_n410_ | ~new_n411_)) | (new_n408_ & (~\a[23]  ^ (new_n407_ & (~new_n98_ | ~new_n406_)))) | (~new_n408_ & (~\a[23]  | ~new_n407_ | (new_n98_ & new_n406_)) & (\a[23]  | (new_n407_ & (~new_n98_ | ~new_n406_)))));
  assign new_n406_ = (\a[20]  | \a[21] ) & (~\a[20]  | ~\a[21] ) & (~\a[22]  | ~\a[23] ) & (\a[22]  | \a[23] );
  assign new_n407_ = (~\b[2]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  ^ ~\a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[3]  | (~\a[20]  ^ ~\a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[4]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  ^ \a[23] ));
  assign new_n408_ = ((\b[0]  & (\a[23]  ^ ~\a[24] ) & (~\a[24]  | ~\a[25] ) & (\a[24]  | \a[25] )) | (\b[1]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] ) & (~\a[25]  ^ \a[26] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] ) & (~\a[25]  | ~\a[26] ) & (\a[25]  | \a[26] ))) ^ (\a[26]  & \b[0]  & (\a[23]  | \a[24] ) & (~\a[23]  | ~\a[24] ));
  assign new_n409_ = \b[0]  & (~\a[23]  | ~\a[24] ) & (\a[23]  | \a[24] ) & (~\b[0]  | (~\a[20]  ^ ~\a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[1]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  ^ \a[23] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] )) & \a[23]  & (~\b[0]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~\b[0]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  ^ ~\a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[1]  | (~\a[20]  ^ ~\a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[2]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  ^ \a[23] )) & ((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )));
  assign new_n410_ = \a[23]  ^ (((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  ^ ~\a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[2]  | (~\a[20]  ^ ~\a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[3]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  ^ \a[23] )));
  assign new_n411_ = (\b[0]  & (~\a[23]  | ~\a[24] ) & (\a[23]  | \a[24] )) ^ ((~\b[0]  | (~\a[20]  ^ ~\a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[1]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  ^ \a[23] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] )) & \a[23]  & (~\b[0]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] )) & (~\b[0]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  ^ ~\a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[1]  | (~\a[20]  ^ ~\a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[2]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  ^ \a[23] )) & ((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n412_ = (~\a[26]  | ((~\b[0]  | (~\a[23]  ^ ~\a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[1]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  ^ \a[26] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )) & \a[26]  & (~\b[0]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] )))) ^ ((~\b[1]  | (~\a[23]  ^ ~\a[24] ) | (\a[24]  & \a[25] ) | (~\a[24]  & ~\a[25] )) & (~\b[2]  | (~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  ^ \a[26] )) & ((~\a[23]  & ~\a[24] ) | (\a[23]  & \a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (\a[24]  ^ \a[25] ) | (~\a[23]  ^ ~\a[24] ) | (\a[25]  & \a[26] ) | (~\a[25]  & ~\a[26] )));
  assign new_n413_ = ~new_n398_ ^ ((new_n303_ ^ ~new_n304_) ^ ((~new_n305_ & new_n313_) | (~new_n306_ & (new_n305_ | ~new_n313_) & (~new_n305_ | new_n313_))));
  assign new_n414_ = \a[23]  ^ (new_n415_ & (~new_n406_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n415_ = (~\b[8]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  ^ ~\a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[9]  | (~\a[20]  ^ ~\a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[10]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  ^ \a[23] ));
  assign new_n416_ = \a[23]  ^ ((~\b[6]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[7]  | (\a[20]  ^ \a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[8]  | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  ^ \a[23] )) & ((\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n79_ & (~\b[7]  ^ \b[8] ))));
  assign new_n417_ = ~new_n393_ ^ (new_n300_ ^ ~new_n392_);
  assign new_n418_ = ~new_n390_ ^ (new_n314_ ^ ((~new_n317_ & (new_n233_ | (~new_n232_ & new_n240_) | (new_n232_ & ~new_n240_)) & (~new_n233_ | (~new_n232_ ^ new_n240_))) | (~new_n300_ & (new_n317_ | (~new_n233_ & (new_n232_ | ~new_n240_) & (~new_n232_ | new_n240_)) | (new_n233_ & (new_n232_ ^ new_n240_))) & (~new_n317_ | (~new_n233_ ^ (~new_n232_ ^ new_n240_))))));
  assign new_n419_ = \a[23]  ^ ((~\b[11]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[12]  | (\a[20]  ^ \a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[13]  | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  ^ \a[23] )) & (~new_n133_ | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] )));
  assign new_n420_ = new_n385_ & (~new_n291_ ^ (new_n292_ | (~new_n295_ & new_n318_)));
  assign new_n421_ = \a[23]  ^ ((~\b[14]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[15]  | (\a[20]  ^ \a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[16]  | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  ^ \a[23] )) & (~new_n186_ | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] )));
  assign new_n422_ = \a[23]  ^ ((~\b[12]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[13]  | (\a[20]  ^ \a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[14]  | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  ^ \a[23] )) & ((\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n142_ & (~\b[13]  ^ \b[14] ))));
  assign new_n423_ = ~new_n381_ ^ (new_n286_ ^ ~new_n380_);
  assign new_n424_ = ~new_n378_ ^ ((~new_n284_ & ~new_n320_) ^ ((~new_n322_ & (new_n222_ | ~new_n282_) & (~new_n222_ | new_n282_)) | (~new_n286_ & (new_n322_ | (~new_n222_ & new_n282_) | (new_n222_ & ~new_n282_)) & (~new_n322_ | (~new_n222_ ^ new_n282_)))));
  assign new_n425_ = \a[23]  ^ ((~\b[17]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[18]  | (\a[20]  ^ \a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[19]  | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  ^ \a[23] )) & (~new_n253_ | (\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] )));
  assign new_n426_ = ~new_n373_ ^ ((~new_n278_ ^ new_n325_) ^ ((~new_n326_ & (~new_n216_ | new_n323_) & (new_n216_ | ~new_n323_)) | (~new_n279_ & (new_n326_ | (new_n216_ & ~new_n323_) | (~new_n216_ & new_n323_)) & (~new_n326_ | (new_n216_ ^ ~new_n323_)))));
  assign new_n427_ = ~new_n326_ ^ (new_n216_ ^ ~new_n323_);
  assign new_n428_ = \a[23]  ^ (((\a[20]  & \a[21] ) | (~\a[20]  & ~\a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~new_n201_ ^ ~\b[19] )) & (~\b[18]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\a[20]  ^ \a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[19]  | (\a[20]  ^ \a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )));
  assign new_n429_ = (~new_n430_ | ~\a[20] ) & ((~new_n430_ & ~\a[20] ) | (new_n430_ & \a[20] ) | ((~\a[20]  | ((~new_n365_ | ~\a[23] ) & (new_n365_ | \a[23] ) & ((new_n367_ & \a[23] ) | ((~new_n367_ | ~\a[23] ) & (new_n367_ | \a[23] ) & ((new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] )))))) | ((~new_n365_ ^ \a[23] ) & (~new_n367_ | ~\a[23] ) & ((new_n367_ & \a[23] ) | (~new_n367_ & ~\a[23] ) | ((~new_n368_ | ~\a[23] ) & (new_n370_ | (new_n368_ & \a[23] ) | (~new_n368_ & ~\a[23] )))))) & (((~\a[20]  | ((~new_n367_ | ~\a[23] ) & (new_n367_ | \a[23] ) & ((new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] )))) | ((~new_n367_ ^ \a[23] ) & (~new_n368_ | ~\a[23] ) & (new_n370_ | (new_n368_ & \a[23] ) | (~new_n368_ & ~\a[23] )))) & (new_n431_ | (\a[20]  & ((new_n367_ & \a[23] ) | (~new_n367_ & ~\a[23] ) | ((~new_n368_ | ~\a[23] ) & (new_n370_ | (new_n368_ & \a[23] ) | (~new_n368_ & ~\a[23] )))) & ((new_n367_ ^ \a[23] ) | (new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] )))) | (~\a[20]  & ((~new_n367_ ^ \a[23] ) ^ ((new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] ))))))) | (\a[20]  & ((new_n365_ & \a[23] ) | (~new_n365_ & ~\a[23] ) | ((~new_n367_ | ~\a[23] ) & ((new_n367_ & \a[23] ) | (~new_n367_ & ~\a[23] ) | ((~new_n368_ | ~\a[23] ) & (new_n370_ | (new_n368_ & \a[23] ) | (~new_n368_ & ~\a[23] )))))) & ((new_n365_ ^ \a[23] ) | (new_n367_ & \a[23] ) | ((~new_n367_ | ~\a[23] ) & (new_n367_ | \a[23] ) & ((new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] )))))) | (~\a[20]  & ((~new_n365_ ^ \a[23] ) ^ ((new_n367_ & \a[23] ) | ((~new_n367_ | ~\a[23] ) & (new_n367_ | \a[23] ) & ((new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] ))))))))));
  assign new_n430_ = ((new_n365_ & \a[23] ) | ((~new_n365_ | ~\a[23] ) & (new_n365_ | \a[23] ) & ((new_n367_ & \a[23] ) | (((new_n368_ & \a[23] ) | (~new_n370_ & (new_n368_ | \a[23] ) & (~new_n368_ | ~\a[23] ))) & (~new_n367_ | ~\a[23] ) & (new_n367_ | \a[23] ))))) ^ (\a[23]  ^ (new_n268_ ^ ~new_n364_));
  assign new_n431_ = (~\a[20]  | (new_n370_ & ~new_n432_) | (~new_n370_ & new_n432_)) & (((~new_n433_ | ~\a[20] ) & ((new_n433_ & \a[20] ) | (~new_n433_ & ~\a[20] ) | ((~new_n434_ | ~\a[20] ) & (((~new_n435_ | ~\a[20] ) & (new_n436_ | (~new_n435_ & ~\a[20] ) | (new_n435_ & \a[20] ))) | (new_n434_ & \a[20] ) | (~new_n434_ & ~\a[20] ))))) | (\a[20]  & (~new_n370_ | new_n432_) & (new_n370_ | ~new_n432_)) | (~\a[20]  & (~new_n370_ ^ ~new_n432_)));
  assign new_n432_ = \a[23]  ^ (new_n275_ ^ ~new_n369_);
  assign new_n433_ = (new_n371_ ^ \a[23] ) ^ (new_n372_ | (new_n426_ & ((~new_n428_ & (new_n279_ | ~new_n427_) & (~new_n279_ | new_n427_)) | (~new_n374_ & (new_n428_ | (~new_n279_ & new_n427_) | (new_n279_ & ~new_n427_)) & (~new_n428_ | (~new_n279_ ^ new_n427_))))));
  assign new_n434_ = new_n426_ ^ ((~new_n428_ & (~new_n279_ | new_n427_) & (new_n279_ | ~new_n427_)) | (~new_n374_ & (new_n428_ | (new_n279_ & ~new_n427_) | (~new_n279_ & new_n427_)) & (~new_n428_ | (new_n279_ ^ ~new_n427_))));
  assign new_n435_ = ~new_n374_ ^ (~new_n428_ ^ (~new_n279_ ^ new_n427_));
  assign new_n436_ = (~new_n437_ | ~\a[20] ) & ((new_n437_ & \a[20] ) | (~new_n437_ & ~\a[20] ) | (~new_n438_ & (new_n438_ | new_n492_ | ((new_n493_ | (~new_n382_ & new_n423_) | (new_n382_ & ~new_n423_)) & (new_n440_ | (~new_n493_ & (new_n382_ | ~new_n423_) & (~new_n382_ | new_n423_)) | (new_n493_ & (new_n382_ ^ new_n423_)))))));
  assign new_n437_ = (new_n375_ ^ ~new_n425_) ^ (new_n377_ | (new_n424_ & (new_n379_ | (~new_n382_ & new_n423_))));
  assign new_n438_ = ~new_n439_ & (~new_n424_ | (~new_n379_ & (new_n382_ | ~new_n423_))) & (new_n424_ | new_n379_ | (~new_n382_ & new_n423_));
  assign new_n439_ = \a[20]  ^ (~\b[19]  | (((\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (new_n201_ | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ))));
  assign new_n440_ = (~new_n441_ | new_n491_) & ((new_n441_ & ~new_n491_) | (~new_n441_ & new_n491_) | (~new_n443_ & (~new_n490_ | (~new_n445_ & (new_n448_ | ~new_n489_)))));
  assign new_n441_ = new_n442_ ^ (new_n384_ | (((~new_n422_ & (new_n295_ | ~new_n318_) & (~new_n295_ | new_n318_)) | (~new_n386_ & (new_n422_ | (~new_n295_ & new_n318_) | (new_n295_ & ~new_n318_)) & (~new_n422_ | (~new_n295_ ^ new_n318_)))) & ~new_n384_ & ~new_n420_));
  assign new_n442_ = ~new_n421_ ^ ((new_n287_ ^ ~new_n319_) ^ (new_n289_ | (new_n291_ & (new_n292_ | (~new_n295_ & new_n318_)))));
  assign new_n443_ = ~new_n444_ & (new_n384_ | new_n420_ | ((new_n422_ | (~new_n295_ & new_n318_) | (new_n295_ & ~new_n318_)) & (new_n386_ | (~new_n422_ & (new_n295_ | ~new_n318_) & (~new_n295_ | new_n318_)) | (new_n422_ & (new_n295_ ^ new_n318_))))) & ((~new_n384_ & ~new_n420_) | (~new_n422_ & (new_n295_ | ~new_n318_) & (~new_n295_ | new_n318_)) | (~new_n386_ & (new_n422_ | (~new_n295_ & new_n318_) | (new_n295_ & ~new_n318_)) & (~new_n422_ | (~new_n295_ ^ new_n318_))));
  assign new_n444_ = \a[20]  ^ ((~\b[16]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[17]  | (\a[17]  ^ \a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[18]  | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  ^ \a[20] )) & (~new_n199_ | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n445_ = ~new_n447_ & (~new_n386_ | new_n446_) & (new_n386_ | ~new_n446_);
  assign new_n446_ = ~new_n422_ ^ (new_n295_ ^ ~new_n318_);
  assign new_n447_ = \a[20]  ^ ((~\b[15]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[16]  | (\a[17]  ^ \a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[17]  | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  ^ \a[20] )) & (~new_n144_ | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n448_ = (~new_n449_ | new_n487_) & ((new_n449_ & ~new_n487_) | (~new_n449_ & new_n487_) | (~new_n450_ & (new_n450_ | new_n486_ | ((new_n488_ | (~new_n394_ & new_n417_) | (new_n394_ & ~new_n417_)) & (new_n452_ | (~new_n488_ & (new_n394_ | ~new_n417_) & (~new_n394_ | new_n417_)) | (new_n488_ & (new_n394_ ^ new_n417_)))))));
  assign new_n449_ = (new_n387_ ^ ~new_n419_) ^ (new_n389_ | (new_n418_ & (new_n391_ | (~new_n394_ & new_n417_))));
  assign new_n450_ = ~new_n451_ & (~new_n418_ | (~new_n391_ & (new_n394_ | ~new_n417_))) & (new_n418_ | new_n391_ | (~new_n394_ & new_n417_));
  assign new_n451_ = \a[20]  ^ ((((~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] ) & ((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )))) | ((~\b[14]  ^ \b[15] ) & (~\b[13]  | ~\b[14] ) & (new_n142_ | (\b[13]  & \b[14] ) | (~\b[13]  & ~\b[14] ))) | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )) & (~\b[13]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[14]  | (\a[17]  ^ \a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[15]  | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  ^ \a[20] )));
  assign new_n452_ = (~new_n453_ | new_n485_) & ((new_n453_ & ~new_n485_) | (~new_n453_ & new_n485_) | (~new_n455_ & (~new_n484_ | (~new_n457_ & (new_n460_ | ~new_n483_)))));
  assign new_n453_ = new_n454_ ^ (new_n397_ | (new_n413_ & ((~new_n416_ & (new_n306_ | (~new_n305_ & new_n313_) | (new_n305_ & ~new_n313_)) & (~new_n306_ | (~new_n305_ ^ new_n313_))) | (~new_n399_ & (new_n416_ | (~new_n306_ & (new_n305_ | ~new_n313_) & (~new_n305_ | new_n313_)) | (new_n306_ & (new_n305_ ^ new_n313_))) & (~new_n416_ | (~new_n306_ ^ (~new_n305_ ^ new_n313_)))))));
  assign new_n454_ = ~new_n414_ ^ ((new_n301_ ^ ~new_n302_) ^ ((new_n303_ & ~new_n304_) | ((~new_n303_ | new_n304_) & (new_n303_ | ~new_n304_) & ((~new_n305_ & new_n313_) | (~new_n306_ & (new_n305_ | ~new_n313_) & (~new_n305_ | new_n313_))))));
  assign new_n455_ = ~new_n456_ & (~new_n413_ | ((new_n416_ | (~new_n306_ & (new_n305_ | ~new_n313_) & (~new_n305_ | new_n313_)) | (new_n306_ & (new_n305_ ^ new_n313_))) & (new_n399_ | (~new_n416_ & (new_n306_ | (~new_n305_ & new_n313_) | (new_n305_ & ~new_n313_)) & (~new_n306_ | (~new_n305_ ^ new_n313_))) | (new_n416_ & (new_n306_ ^ (~new_n305_ ^ new_n313_)))))) & (new_n413_ | (~new_n416_ & (new_n306_ | (~new_n305_ & new_n313_) | (new_n305_ & ~new_n313_)) & (~new_n306_ | (~new_n305_ ^ new_n313_))) | (~new_n399_ & (new_n416_ | (~new_n306_ & (new_n305_ | ~new_n313_) & (~new_n305_ | new_n313_)) | (new_n306_ & (new_n305_ ^ new_n313_))) & (~new_n416_ | (~new_n306_ ^ (~new_n305_ ^ new_n313_)))));
  assign new_n456_ = \a[20]  ^ ((~\b[10]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[11]  | (\a[17]  ^ \a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[12]  | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  ^ \a[20] )) & (~new_n107_ | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n457_ = ~new_n459_ & (~new_n399_ | new_n458_) & (new_n399_ | ~new_n458_);
  assign new_n458_ = ~new_n416_ ^ (~new_n306_ ^ (~new_n305_ ^ new_n313_));
  assign new_n459_ = \a[20]  ^ ((~\b[9]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[10]  | (\a[17]  ^ \a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[11]  | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  ^ \a[20] )) & (~new_n135_ | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n460_ = (~new_n462_ | new_n480_) & ((~new_n463_ & (~new_n479_ | ((new_n482_ | (new_n461_ & ~new_n405_) | (~new_n461_ & new_n405_)) & (new_n465_ | (~new_n482_ & (~new_n461_ | new_n405_) & (new_n461_ | ~new_n405_)) | (new_n482_ & (~new_n461_ ^ ~new_n405_)))))) | (new_n462_ & ~new_n480_) | (~new_n462_ & new_n480_));
  assign new_n461_ = new_n404_ ^ ~new_n412_;
  assign new_n462_ = (new_n400_ ^ ~new_n401_) ^ ((new_n402_ & ~new_n403_) | (((~new_n404_ & new_n412_) | (~new_n405_ & (new_n404_ | ~new_n412_) & (~new_n404_ | new_n412_))) & (~new_n402_ | new_n403_) & (new_n402_ | ~new_n403_)));
  assign new_n463_ = ~new_n464_ & ((new_n402_ & ~new_n403_) | (~new_n402_ & new_n403_) | ((new_n404_ | ~new_n412_) & (new_n405_ | (~new_n404_ & new_n412_) | (new_n404_ & ~new_n412_)))) & ((new_n402_ ^ ~new_n403_) | (~new_n404_ & new_n412_) | (~new_n405_ & (new_n404_ | ~new_n412_) & (~new_n404_ | new_n412_)));
  assign new_n464_ = \a[20]  ^ ((((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))) | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )) & (~\b[7]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[8]  | (\a[17]  ^ \a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[9]  | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  ^ \a[20] )));
  assign new_n465_ = (new_n466_ | ~new_n467_) & ((new_n466_ & ~new_n467_) | (~new_n466_ & new_n467_) | ((~new_n468_ | new_n469_) & (((new_n470_ | ~new_n478_) & (new_n471_ | (~new_n470_ & new_n478_) | (new_n470_ & ~new_n478_))) | (new_n468_ & ~new_n469_) | (~new_n468_ & new_n469_))));
  assign new_n466_ = \a[20]  ^ ((~\b[5]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[6]  | (\a[17]  ^ \a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[7]  | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  ^ \a[20] )) & (~new_n88_ | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n467_ = (new_n409_ | (~new_n410_ & new_n411_)) ^ (new_n408_ ^ (~\a[23]  ^ (new_n407_ & (~new_n98_ | ~new_n406_))));
  assign new_n468_ = new_n410_ ^ ~new_n411_;
  assign new_n469_ = \a[20]  ^ ((~\b[4]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[5]  | (\a[17]  ^ \a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[6]  | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  ^ \a[20] )) & (~new_n91_ | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n470_ = \a[20]  ^ ((~\b[3]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[4]  | (\a[17]  ^ \a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[5]  | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  ^ \a[20] )) & (~new_n94_ | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n471_ = (~new_n474_ | (\a[20]  ^ (new_n473_ & (~new_n98_ | ~new_n472_)))) & ((~new_n475_ & (new_n476_ | ~new_n477_)) | (new_n474_ & (~\a[20]  ^ (new_n473_ & (~new_n98_ | ~new_n472_)))) | (~new_n474_ & (~\a[20]  | ~new_n473_ | (new_n98_ & new_n472_)) & (\a[20]  | (new_n473_ & (~new_n98_ | ~new_n472_)))));
  assign new_n472_ = (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ) & (~\a[19]  | ~\a[20] ) & (\a[19]  | \a[20] );
  assign new_n473_ = (~\b[2]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  ^ ~\a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[3]  | (~\a[17]  ^ ~\a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[4]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  ^ \a[20] ));
  assign new_n474_ = ((\b[0]  & (\a[20]  ^ ~\a[21] ) & (~\a[21]  | ~\a[22] ) & (\a[21]  | \a[22] )) | (\b[1]  & (\a[20]  | \a[21] ) & (~\a[20]  | ~\a[21] ) & (~\a[22]  ^ \a[23] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & (\a[20]  | \a[21] ) & (~\a[20]  | ~\a[21] ) & (~\a[22]  | ~\a[23] ) & (\a[22]  | \a[23] ))) ^ (\a[23]  & \b[0]  & (\a[20]  | \a[21] ) & (~\a[20]  | ~\a[21] ));
  assign new_n475_ = \b[0]  & (~\a[20]  | ~\a[21] ) & (\a[20]  | \a[21] ) & (~\b[0]  | (~\a[17]  ^ ~\a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[1]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  ^ \a[20] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )) & \a[20]  & (~\b[0]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[0]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  ^ ~\a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[1]  | (~\a[17]  ^ ~\a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[2]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  ^ \a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )));
  assign new_n476_ = \a[20]  ^ (((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  ^ ~\a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[2]  | (~\a[17]  ^ ~\a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[3]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  ^ \a[20] )));
  assign new_n477_ = (\b[0]  & (~\a[20]  | ~\a[21] ) & (\a[20]  | \a[21] )) ^ ((~\b[0]  | (~\a[17]  ^ ~\a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[1]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  ^ \a[20] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )) & \a[20]  & (~\b[0]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[0]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  ^ ~\a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[1]  | (~\a[17]  ^ ~\a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[2]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  ^ \a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n478_ = ((~\b[0]  | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (~\a[20]  ^ ~\a[21] ) | (\a[21]  ^ \a[22] )) & (~\b[1]  | (~\a[20]  ^ ~\a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[2]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  ^ \a[23] )) & ((~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))) ^ (~\a[23]  | ((~\b[0]  | (~\a[20]  ^ ~\a[21] ) | (\a[21]  & \a[22] ) | (~\a[21]  & ~\a[22] )) & (~\b[1]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  ^ \a[23] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ) | (\a[22]  & \a[23] ) | (~\a[22]  & ~\a[23] )) & \a[23]  & (~\b[0]  | (~\a[20]  & ~\a[21] ) | (\a[20]  & \a[21] ))));
  assign new_n479_ = ~new_n464_ ^ ((new_n402_ ^ ~new_n403_) ^ ((~new_n404_ & new_n412_) | (~new_n405_ & (new_n404_ | ~new_n412_) & (~new_n404_ | new_n412_))));
  assign new_n480_ = \a[20]  ^ (new_n481_ & (~new_n472_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n481_ = (~\b[8]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  ^ ~\a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[9]  | (~\a[17]  ^ ~\a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[10]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  ^ \a[20] ));
  assign new_n482_ = \a[20]  ^ ((~\b[6]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[7]  | (\a[17]  ^ \a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[8]  | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  ^ \a[20] )) & ((\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n79_ & (~\b[7]  ^ \b[8] ))));
  assign new_n483_ = ~new_n459_ ^ (new_n399_ ^ ~new_n458_);
  assign new_n484_ = ~new_n456_ ^ (new_n413_ ^ ((~new_n416_ & (new_n306_ | (~new_n305_ & new_n313_) | (new_n305_ & ~new_n313_)) & (~new_n306_ | (~new_n305_ ^ new_n313_))) | (~new_n399_ & (new_n416_ | (~new_n306_ & (new_n305_ | ~new_n313_) & (~new_n305_ | new_n313_)) | (new_n306_ & (new_n305_ ^ new_n313_))) & (~new_n416_ | (~new_n306_ ^ (~new_n305_ ^ new_n313_))))));
  assign new_n485_ = \a[20]  ^ ((~\b[11]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[12]  | (\a[17]  ^ \a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[13]  | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  ^ \a[20] )) & (~new_n133_ | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n486_ = new_n451_ & (~new_n418_ ^ (new_n391_ | (~new_n394_ & new_n417_)));
  assign new_n487_ = \a[20]  ^ ((~\b[14]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[15]  | (\a[17]  ^ \a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[16]  | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  ^ \a[20] )) & (~new_n186_ | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n488_ = \a[20]  ^ ((~\b[12]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[13]  | (\a[17]  ^ \a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[14]  | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  ^ \a[20] )) & ((\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n142_ & (~\b[13]  ^ \b[14] ))));
  assign new_n489_ = ~new_n447_ ^ (new_n386_ ^ ~new_n446_);
  assign new_n490_ = ~new_n444_ ^ ((~new_n384_ & ~new_n420_) ^ ((~new_n422_ & (new_n295_ | ~new_n318_) & (~new_n295_ | new_n318_)) | (~new_n386_ & (new_n422_ | (~new_n295_ & new_n318_) | (new_n295_ & ~new_n318_)) & (~new_n422_ | (~new_n295_ ^ new_n318_)))));
  assign new_n491_ = \a[20]  ^ ((~\b[17]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[18]  | (\a[17]  ^ \a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[19]  | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  ^ \a[20] )) & (~new_n253_ | (\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )));
  assign new_n492_ = new_n439_ & (~new_n424_ ^ (new_n379_ | (~new_n382_ & new_n423_)));
  assign new_n493_ = \a[20]  ^ (((\a[17]  & \a[18] ) | (~\a[17]  & ~\a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~new_n201_ ^ ~\b[19] )) & (~\b[18]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\a[17]  ^ \a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[19]  | (\a[17]  ^ \a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )));
  assign new_n494_ = ((new_n508_ & \a[23] ) | ((new_n508_ | \a[23] ) & (~new_n508_ | ~\a[23] ) & ((new_n495_ & \a[23] ) | (~new_n507_ & (~new_n495_ | ~\a[23] ) & (new_n495_ | \a[23] ))))) ^ (\a[23]  ^ (~new_n520_ ^ (~new_n521_ ^ ~\a[26] )));
  assign new_n495_ = (new_n496_ ^ \a[26] ) ^ ((\a[26]  & ((new_n347_ & \a[29] ) | (~new_n347_ & ~\a[29] ) | ((~new_n334_ | ~\a[29] ) & (new_n331_ | (~new_n334_ & ~\a[29] ) | (new_n334_ & \a[29] )))) & ((new_n347_ ^ \a[29] ) | (new_n334_ & \a[29] ) | (~new_n331_ & (new_n334_ | \a[29] ) & (~new_n334_ | ~\a[29] )))) | (~new_n345_ & (~\a[26]  | ((~new_n347_ | ~\a[29] ) & (new_n347_ | \a[29] ) & ((new_n334_ & \a[29] ) | (~new_n331_ & (new_n334_ | \a[29] ) & (~new_n334_ | ~\a[29] )))) | ((~new_n347_ ^ \a[29] ) & (~new_n334_ | ~\a[29] ) & (new_n331_ | (~new_n334_ & ~\a[29] ) | (new_n334_ & \a[29] )))) & (\a[26]  | ((new_n347_ ^ \a[29] ) ^ ((new_n334_ & \a[29] ) | (~new_n331_ & (new_n334_ | \a[29] ) & (~new_n334_ | ~\a[29] )))))));
  assign new_n496_ = (new_n497_ ^ \a[29] ) ^ ((new_n347_ & \a[29] ) | ((new_n347_ | \a[29] ) & (~new_n347_ | ~\a[29] ) & ((new_n334_ & \a[29] ) | (~new_n331_ & (~new_n334_ | ~\a[29] ) & (new_n334_ | \a[29] )))));
  assign new_n497_ = (~new_n498_ & (~new_n349_ | (~new_n348_ & ~new_n360_))) ^ (~new_n499_ ^ \a[32] );
  assign new_n498_ = ~new_n359_ & (~new_n350_ | new_n352_) & (new_n350_ | ~new_n352_);
  assign new_n499_ = new_n501_ ^ (new_n500_ | (~new_n350_ & new_n352_));
  assign new_n500_ = ~new_n354_ & (~new_n355_ | (~new_n358_ & (new_n353_ | ~new_n340_))) & (new_n355_ | new_n358_ | (~new_n353_ & new_n340_));
  assign new_n501_ = ~new_n506_ ^ (new_n503_ ^ (new_n502_ | new_n505_));
  assign new_n502_ = new_n355_ & (new_n358_ | (new_n340_ & (new_n342_ | (new_n261_ & (new_n263_ | (new_n192_ & ~new_n194_))))));
  assign new_n503_ = ~new_n504_ ^ (\a[38]  & ~\b[13] );
  assign new_n504_ = (~\b[14]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (\a[35]  ^ \a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[15]  | (\a[35]  ^ \a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[16]  | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  ^ \a[38] )) & (~new_n186_ | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ));
  assign new_n505_ = \a[38]  & \b[12]  & new_n357_ & (~new_n356_ | ~new_n80_);
  assign new_n506_ = \a[35]  ^ ((~new_n253_ | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & (~\b[18]  | (\a[32]  ^ \a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[19]  | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  ^ \a[35] )) & (~\b[17]  | (\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )));
  assign new_n507_ = (~\a[23]  | (new_n345_ & ~new_n346_) | (~new_n345_ & new_n346_)) & (((~\a[23]  | (new_n71_ & ~new_n330_) | (~new_n71_ & new_n330_)) & ((\a[23]  & (~new_n71_ | new_n330_) & (new_n71_ | ~new_n330_)) | (~\a[23]  & (~new_n71_ ^ ~new_n330_)) | ((~new_n361_ | ~\a[23] ) & ((new_n361_ & \a[23] ) | (~new_n361_ & ~\a[23] ) | ((~new_n362_ | ~\a[23] ) & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] ))))))) | (\a[23]  & (~new_n345_ | new_n346_) & (new_n345_ | ~new_n346_)) | (~\a[23]  & (~new_n345_ ^ ~new_n346_)));
  assign new_n508_ = (new_n510_ ^ \a[26] ) ^ ((new_n496_ & \a[26] ) | ((~new_n496_ | ~\a[26] ) & (new_n496_ | \a[26] ) & ((\a[26]  & (~new_n509_ | (~new_n519_ & (new_n331_ | ~new_n333_))) & (new_n509_ | new_n519_ | (~new_n331_ & new_n333_))) | (((\a[26]  & (new_n331_ | ~new_n333_) & (~new_n331_ | new_n333_)) | (~new_n71_ & (~\a[26]  | (~new_n331_ & new_n333_) | (new_n331_ & ~new_n333_)) & (\a[26]  | (~new_n331_ ^ new_n333_)))) & (~\a[26]  | (new_n509_ & (new_n519_ | (~new_n331_ & new_n333_))) | (~new_n509_ & ~new_n519_ & (new_n331_ | ~new_n333_))) & (\a[26]  | (new_n509_ ^ (new_n519_ | (~new_n331_ & new_n333_))))))));
  assign new_n509_ = ~new_n347_ ^ ~\a[29] ;
  assign new_n510_ = (new_n511_ ^ \a[29] ) ^ ((new_n497_ & \a[29] ) | ((new_n497_ | \a[29] ) & (~new_n497_ | ~\a[29] ) & ((new_n347_ & \a[29] ) | ((~new_n347_ | ~\a[29] ) & (new_n347_ | \a[29] ) & ((new_n334_ & \a[29] ) | (~new_n331_ & (~new_n334_ | ~\a[29] ) & (new_n334_ | \a[29] )))))));
  assign new_n511_ = (~new_n512_ ^ ~\a[32] ) ^ ((new_n499_ & \a[32] ) | ((~new_n499_ | ~\a[32] ) & (new_n499_ | \a[32] ) & (new_n498_ | (new_n349_ & (new_n348_ | new_n360_)))));
  assign new_n512_ = new_n514_ ^ ((new_n513_ & ~new_n506_) | (new_n501_ & (new_n500_ | (~new_n350_ & new_n352_))));
  assign new_n513_ = new_n503_ ^ (new_n502_ | new_n505_);
  assign new_n514_ = ~new_n518_ ^ (new_n515_ ^ (new_n517_ | (new_n503_ & (new_n502_ | new_n505_))));
  assign new_n515_ = ~new_n516_ ^ (\a[38]  & ~\b[14] );
  assign new_n516_ = (~\b[15]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (\a[35]  ^ \a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[16]  | (\a[35]  ^ \a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[17]  | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  ^ \a[38] )) & (~new_n144_ | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ));
  assign new_n517_ = new_n504_ & \a[38]  & \b[13] ;
  assign new_n518_ = \a[35]  ^ (((\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] ) | (~new_n201_ ^ ~\b[19] )) & (~\b[19]  | (\a[32]  ^ \a[33] ) | (\a[33]  & \a[34] ) | (~\a[33]  & ~\a[34] )) & (~\b[18]  | (\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )));
  assign new_n519_ = new_n334_ & \a[29] ;
  assign new_n520_ = (~new_n510_ | ~\a[26] ) & ((new_n510_ & \a[26] ) | (~new_n510_ & ~\a[26] ) | ((~new_n496_ | ~\a[26] ) & ((new_n496_ & \a[26] ) | (~new_n496_ & ~\a[26] ) | ((~\a[26]  | (new_n509_ & (new_n519_ | (~new_n331_ & new_n333_))) | (~new_n509_ & ~new_n519_ & (new_n331_ | ~new_n333_))) & (((~\a[26]  | (~new_n331_ & new_n333_) | (new_n331_ & ~new_n333_)) & (new_n71_ | (\a[26]  & (new_n331_ | ~new_n333_) & (~new_n331_ | new_n333_)) | (~\a[26]  & (new_n331_ ^ new_n333_)))) | (\a[26]  & (~new_n509_ | (~new_n519_ & (new_n331_ | ~new_n333_))) & (new_n509_ | new_n519_ | (~new_n331_ & new_n333_))) | (~\a[26]  & (~new_n509_ ^ (new_n519_ | (~new_n331_ & new_n333_)))))))));
  assign new_n521_ = ((new_n511_ & \a[29] ) | ((~new_n511_ | ~\a[29] ) & (new_n511_ | \a[29] ) & ((new_n497_ & \a[29] ) | ((~new_n497_ | ~\a[29] ) & (new_n497_ | \a[29] ) & ((new_n347_ & \a[29] ) | (((new_n334_ & \a[29] ) | (~new_n331_ & (~new_n334_ | ~\a[29] ) & (new_n334_ | \a[29] ))) & (~new_n347_ | ~\a[29] ) & (new_n347_ | \a[29] ))))))) ^ (\a[29]  ^ (~new_n522_ ^ new_n523_));
  assign new_n522_ = (~new_n512_ | ~\a[32] ) & ((~new_n512_ & ~\a[32] ) | (new_n512_ & \a[32] ) | ((~new_n499_ | ~\a[32] ) & ((new_n499_ & \a[32] ) | (~new_n499_ & ~\a[32] ) | (~new_n498_ & (~new_n349_ | (~new_n348_ & ~new_n360_))))));
  assign new_n523_ = ~new_n524_ ^ ~\a[32] ;
  assign new_n524_ = new_n526_ ^ (new_n525_ | (new_n514_ & ((new_n513_ & ~new_n506_) | ((new_n513_ | ~new_n506_) & (~new_n513_ | new_n506_) & (new_n500_ | (~new_n350_ & new_n352_))))));
  assign new_n525_ = ~new_n518_ & (~new_n515_ | (~new_n517_ & (~new_n503_ | (~new_n502_ & ~new_n505_)))) & (new_n515_ | new_n517_ | (new_n503_ & (new_n502_ | new_n505_)));
  assign new_n526_ = ~new_n530_ ^ (new_n527_ ^ (new_n529_ | (new_n515_ & (new_n517_ | (new_n503_ & (new_n502_ | new_n505_))))));
  assign new_n527_ = ~new_n528_ ^ (\a[38]  & ~\b[15] );
  assign new_n528_ = (~\b[16]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (\a[35]  ^ \a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[17]  | (\a[35]  ^ \a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[18]  | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  ^ \a[38] )) & (~new_n199_ | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ));
  assign new_n529_ = new_n516_ & \a[38]  & \b[14] ;
  assign new_n530_ = \a[35]  ^ (~\b[19]  | (((\a[33]  ^ \a[34] ) | (\a[32]  ^ \a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] )) & (new_n201_ | (\a[32]  & \a[33] ) | (~\a[32]  & ~\a[33] ) | (\a[34]  & \a[35] ) | (~\a[34]  & ~\a[35] ))));
  assign new_n531_ = ((~\a[23]  | (~new_n520_ & (~new_n521_ | ~\a[26] ) & (new_n521_ | \a[26] )) | (new_n520_ & (~new_n521_ ^ \a[26] ))) & (((~new_n508_ | ~\a[23] ) & ((new_n508_ & \a[23] ) | (~new_n508_ & ~\a[23] ) | ((~new_n495_ | ~\a[23] ) & (new_n507_ | (~new_n495_ & ~\a[23] ) | (new_n495_ & \a[23] ))))) | (\a[23]  & (new_n520_ | (new_n521_ & \a[26] ) | (~new_n521_ & ~\a[26] )) & (~new_n520_ | (new_n521_ ^ \a[26] ))) | (~\a[23]  & (new_n520_ ^ (new_n521_ ^ \a[26] ))))) ^ (~\a[23]  ^ ((~new_n532_ ^ \a[26] ) ^ ((~new_n521_ | ~\a[26] ) & (new_n520_ | (new_n521_ & \a[26] ) | (~new_n521_ & ~\a[26] )))));
  assign new_n532_ = new_n533_ ^ (~\a[29]  ^ (new_n534_ ^ (~new_n535_ ^ \a[32] )));
  assign new_n533_ = (~\a[29]  | (~new_n522_ & new_n523_) | (new_n522_ & ~new_n523_)) & (((~new_n511_ | ~\a[29] ) & ((new_n511_ & \a[29] ) | (~new_n511_ & ~\a[29] ) | ((~new_n497_ | ~\a[29] ) & ((new_n497_ & \a[29] ) | (~new_n497_ & ~\a[29] ) | ((~new_n347_ | ~\a[29] ) & (((~new_n334_ | ~\a[29] ) & (new_n331_ | (new_n334_ & \a[29] ) | (~new_n334_ & ~\a[29] ))) | (new_n347_ & \a[29] ) | (~new_n347_ & ~\a[29] ))))))) | (\a[29]  & (new_n522_ | ~new_n523_) & (~new_n522_ | new_n523_)) | (~\a[29]  & (new_n522_ ^ new_n523_)));
  assign new_n534_ = (~new_n524_ | ~\a[32] ) & (new_n522_ | (new_n524_ & \a[32] ) | (~new_n524_ & ~\a[32] ));
  assign new_n535_ = new_n539_ ^ (new_n536_ | new_n543_);
  assign new_n536_ = ~new_n537_ & new_n526_;
  assign new_n537_ = (new_n518_ | (~new_n538_ & new_n515_) | (new_n538_ & ~new_n515_)) & ((~new_n518_ & (new_n538_ | ~new_n515_) & (~new_n538_ | new_n515_)) | (new_n518_ & (new_n538_ ^ new_n515_)) | ((~new_n513_ | new_n506_) & ((~new_n513_ & new_n506_) | (new_n513_ & ~new_n506_) | (~new_n500_ & (new_n350_ | ~new_n352_)))));
  assign new_n538_ = ~new_n517_ & (~new_n503_ | (~new_n502_ & ~new_n505_));
  assign new_n539_ = ~new_n540_ ^ ~\a[35] ;
  assign new_n540_ = new_n541_ ^ (((new_n528_ | ~\a[38]  | \b[15] ) & (~new_n528_ | (\a[38]  & ~\b[15] )) & ((~new_n538_ & (new_n516_ | ~\a[38]  | \b[14] ) & (~new_n516_ | (\a[38]  & ~\b[14] ))) | (new_n516_ & \a[38]  & \b[14] ))) | (new_n528_ & \a[38]  & \b[15] ));
  assign new_n541_ = ~new_n542_ ^ (\a[38]  & ~\b[16] );
  assign new_n542_ = (~\b[17]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (\a[35]  ^ \a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[18]  | (\a[35]  ^ \a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] )) & (~\b[19]  | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  ^ \a[38] )) & (~new_n253_ | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ));
  assign new_n543_ = ~new_n530_ & (~new_n527_ | (~new_n529_ & (new_n538_ | ~new_n515_))) & (new_n527_ | new_n529_ | (~new_n538_ & new_n515_));
  assign new_n544_ = ((~new_n559_ | ~\a[23] ) & (new_n558_ | (new_n559_ & \a[23] ) | (~new_n559_ & ~\a[23] ))) ^ (new_n545_ ^ ~\a[23] );
  assign new_n545_ = (new_n546_ ^ \a[26] ) ^ ((new_n557_ & \a[26] ) | ((~new_n557_ | ~\a[26] ) & (new_n557_ | \a[26] ) & ((new_n532_ & \a[26] ) | ((new_n532_ | \a[26] ) & (~new_n532_ | ~\a[26] ) & ((new_n521_ & \a[26] ) | (~new_n520_ & (~new_n521_ | ~\a[26] ) & (new_n521_ | \a[26] )))))));
  assign new_n546_ = ((\a[29]  & (~new_n556_ | ((~new_n535_ | ~\a[32] ) & (new_n534_ | (new_n535_ & \a[32] ) | (~new_n535_ & ~\a[32] )))) & (new_n556_ | (new_n535_ & \a[32] ) | (~new_n534_ & (~new_n535_ | ~\a[32] ) & (new_n535_ | \a[32] )))) | (((\a[29]  & (new_n534_ | (new_n535_ & \a[32] ) | (~new_n535_ & ~\a[32] )) & (~new_n534_ | (new_n535_ ^ \a[32] ))) | (~new_n533_ & (~\a[29]  | (~new_n534_ & (~new_n535_ | ~\a[32] ) & (new_n535_ | \a[32] )) | (new_n534_ & (~new_n535_ ^ \a[32] ))) & (\a[29]  | (~new_n534_ ^ (new_n535_ ^ \a[32] ))))) & (~\a[29]  | (new_n556_ & ((new_n535_ & \a[32] ) | (~new_n534_ & (~new_n535_ | ~\a[32] ) & (new_n535_ | \a[32] )))) | (~new_n556_ & (~new_n535_ | ~\a[32] ) & (new_n534_ | (new_n535_ & \a[32] ) | (~new_n535_ & ~\a[32] )))) & (\a[29]  | (new_n556_ ^ ((new_n535_ & \a[32] ) | (~new_n534_ & (~new_n535_ | ~\a[32] ) & (new_n535_ | \a[32] ))))))) ^ (\a[29]  ^ ((new_n552_ ^ \a[32] ) ^ (new_n547_ | (new_n556_ & ((new_n535_ & \a[32] ) | (~new_n534_ & (~new_n535_ | ~\a[32] ) & (new_n535_ | \a[32] )))))));
  assign new_n547_ = \a[32]  & (((~new_n540_ | ~\a[35] ) & (new_n548_ | (new_n540_ & \a[35] ) | (~new_n540_ & ~\a[35] ))) | (~new_n549_ & ~\a[35] ) | (new_n549_ & \a[35] )) & ((new_n540_ & \a[35] ) | (~new_n548_ & (~new_n540_ | ~\a[35] ) & (new_n540_ | \a[35] )) | (~new_n549_ ^ ~\a[35] ));
  assign new_n548_ = ~new_n536_ & ~new_n543_;
  assign new_n549_ = new_n550_ ^ ~new_n551_;
  assign new_n550_ = ((~new_n542_ & \a[38]  & ~\b[16] ) | (new_n542_ & (~\a[38]  | \b[16] )) | (((~new_n528_ & \a[38]  & ~\b[15] ) | (new_n528_ & (~\a[38]  | \b[15] )) | ((new_n538_ | (~new_n516_ & \a[38]  & ~\b[14] ) | (new_n516_ & (~\a[38]  | \b[14] ))) & (~new_n516_ | ~\a[38]  | ~\b[14] ))) & (~new_n528_ | ~\a[38]  | ~\b[15] ))) & (~new_n542_ | ~\a[38]  | ~\b[16] );
  assign new_n551_ = (\a[38]  & ~\b[17] ) ^ (((~new_n201_ ^ \b[19] ) & (~\a[35]  | ~\a[36] ) & (\a[35]  | \a[36] ) & (~\a[37]  | ~\a[38] ) & (\a[37]  | \a[38] )) | (\b[18]  & (~\a[37]  | ~\a[38] ) & (\a[37]  | \a[38] ) & (~\a[35]  ^ \a[36] ) & (~\a[36]  ^ \a[37] )) | (\b[19]  & (~\a[35]  ^ \a[36] ) & (~\a[36]  | ~\a[37] ) & (\a[36]  | \a[37] )));
  assign new_n552_ = ((~new_n549_ | ~\a[35] ) & ((new_n549_ & \a[35] ) | (~new_n549_ & ~\a[35] ) | ((~new_n540_ | ~\a[35] ) & (new_n548_ | (new_n540_ & \a[35] ) | (~new_n540_ & ~\a[35] ))))) ^ (~\a[35]  ^ (new_n553_ ^ new_n555_));
  assign new_n553_ = ~new_n554_ & (new_n550_ | ~new_n551_);
  assign new_n554_ = \a[38]  & \b[17]  & ((new_n201_ ^ \b[19] ) | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] )) & (~\b[18]  | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (\a[35]  ^ \a[36] ) | (\a[36]  ^ \a[37] )) & (~\b[19]  | (\a[35]  ^ \a[36] ) | (\a[36]  & \a[37] ) | (~\a[36]  & ~\a[37] ));
  assign new_n555_ = (\a[38]  & ~\b[18] ) ^ (~\b[19]  | (((\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (\a[35]  ^ \a[36] ) | (\a[36]  ^ \a[37] )) & (new_n201_ | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] ) | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ))));
  assign new_n556_ = \a[32]  ^ ((~new_n549_ ^ \a[35] ) ^ ((~new_n540_ | ~\a[35] ) & ((~new_n536_ & ~new_n543_) | (new_n540_ & \a[35] ) | (~new_n540_ & ~\a[35] ))));
  assign new_n557_ = ((\a[29]  & (~new_n534_ | (~new_n535_ ^ ~\a[32] )) & (new_n534_ | (~new_n535_ & ~\a[32] ) | (new_n535_ & \a[32] ))) | (~new_n533_ & (~\a[29]  | (new_n534_ & (new_n535_ ^ ~\a[32] )) | (~new_n534_ & (new_n535_ | \a[32] ) & (~new_n535_ | ~\a[32] ))) & (\a[29]  | (new_n534_ ^ (new_n535_ ^ ~\a[32] ))))) ^ (~\a[29]  ^ (~new_n556_ ^ ((new_n535_ & \a[32] ) | (~new_n534_ & (new_n535_ | \a[32] ) & (~new_n535_ | ~\a[32] )))));
  assign new_n558_ = (~\a[23]  | ((~new_n532_ ^ \a[26] ) & (~new_n521_ | ~\a[26] ) & (new_n520_ | (new_n521_ & \a[26] ) | (~new_n521_ & ~\a[26] ))) | ((~new_n532_ | ~\a[26] ) & (new_n532_ | \a[26] ) & ((new_n521_ & \a[26] ) | (~new_n520_ & (~new_n521_ | ~\a[26] ) & (new_n521_ | \a[26] ))))) & (((~\a[23]  | (~new_n520_ & (~new_n521_ | ~\a[26] ) & (new_n521_ | \a[26] )) | (new_n520_ & (~new_n521_ ^ \a[26] ))) & (((~new_n508_ | ~\a[23] ) & ((new_n508_ & \a[23] ) | (~new_n508_ & ~\a[23] ) | ((~new_n495_ | ~\a[23] ) & (new_n507_ | (~new_n495_ & ~\a[23] ) | (new_n495_ & \a[23] ))))) | (\a[23]  & (new_n520_ | (new_n521_ & \a[26] ) | (~new_n521_ & ~\a[26] )) & (~new_n520_ | (new_n521_ ^ \a[26] ))) | (~\a[23]  & (new_n520_ ^ (new_n521_ ^ \a[26] ))))) | (\a[23]  & ((new_n532_ ^ \a[26] ) | (new_n521_ & \a[26] ) | (~new_n520_ & (~new_n521_ | ~\a[26] ) & (new_n521_ | \a[26] ))) & ((new_n532_ & \a[26] ) | (~new_n532_ & ~\a[26] ) | ((~new_n521_ | ~\a[26] ) & (new_n520_ | (new_n521_ & \a[26] ) | (~new_n521_ & ~\a[26] ))))) | (~\a[23]  & ((new_n532_ ^ \a[26] ) ^ ((~new_n521_ | ~\a[26] ) & (new_n520_ | (new_n521_ & \a[26] ) | (~new_n521_ & ~\a[26] ))))));
  assign new_n559_ = (new_n557_ ^ \a[26] ) ^ ((new_n532_ & \a[26] ) | ((new_n532_ | \a[26] ) & (~new_n532_ | ~\a[26] ) & ((new_n521_ & \a[26] ) | (~new_n520_ & (~new_n521_ | ~\a[26] ) & (new_n521_ | \a[26] )))));
  assign new_n560_ = ~new_n558_ ^ (new_n559_ ^ \a[23] );
  assign new_n561_ = (~\a[17]  | ((~new_n560_ ^ \a[20] ) & (~new_n531_ | ~\a[20] ) & (new_n68_ | (new_n531_ & \a[20] ) | (~new_n531_ & ~\a[20] ))) | ((~new_n560_ | ~\a[20] ) & (new_n560_ | \a[20] ) & ((new_n531_ & \a[20] ) | (~new_n68_ & (~new_n531_ | ~\a[20] ) & (new_n531_ | \a[20] ))))) & ((\a[17]  & ((new_n560_ ^ \a[20] ) | (new_n531_ & \a[20] ) | (~new_n68_ & (~new_n531_ | ~\a[20] ) & (new_n531_ | \a[20] ))) & ((new_n560_ & \a[20] ) | (~new_n560_ & ~\a[20] ) | ((~new_n531_ | ~\a[20] ) & (new_n68_ | (new_n531_ & \a[20] ) | (~new_n531_ & ~\a[20] ))))) | (~\a[17]  & ((new_n560_ ^ \a[20] ) ^ ((~new_n531_ | ~\a[20] ) & (new_n68_ | (new_n531_ & \a[20] ) | (~new_n531_ & ~\a[20] ))))) | ((~\a[17]  | (~new_n68_ & (~new_n531_ | ~\a[20] ) & (new_n531_ | \a[20] )) | (new_n68_ & (~new_n531_ ^ \a[20] ))) & ((\a[17]  & (new_n68_ | (new_n531_ & \a[20] ) | (~new_n531_ & ~\a[20] )) & (~new_n68_ | (new_n531_ ^ \a[20] ))) | (~\a[17]  & (new_n68_ ^ (new_n531_ ^ \a[20] ))) | ((~new_n562_ | ~\a[17] ) & ((~new_n562_ & ~\a[17] ) | (new_n562_ & \a[17] ) | ((~new_n563_ | ~\a[17] ) & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] ))))))));
  assign new_n562_ = (new_n494_ ^ \a[20] ) ^ ((\a[20]  & ((~new_n508_ & ~\a[23] ) | (new_n508_ & \a[23] ) | ((~new_n495_ | ~\a[23] ) & (new_n507_ | (new_n495_ & \a[23] ) | (~new_n495_ & ~\a[23] )))) & ((~new_n508_ ^ ~\a[23] ) | (new_n495_ & \a[23] ) | (~new_n507_ & (~new_n495_ | ~\a[23] ) & (new_n495_ | \a[23] )))) | (((\a[20]  & (new_n507_ | (new_n495_ & \a[23] ) | (~new_n495_ & ~\a[23] )) & (~new_n507_ | (new_n495_ ^ \a[23] ))) | (~new_n69_ & (~\a[20]  | (~new_n507_ & (~new_n495_ | ~\a[23] ) & (new_n495_ | \a[23] )) | (new_n507_ & (~new_n495_ ^ \a[23] ))) & (\a[20]  | (~new_n507_ ^ (new_n495_ ^ \a[23] ))))) & (~\a[20]  | ((new_n508_ | \a[23] ) & (~new_n508_ | ~\a[23] ) & ((new_n495_ & \a[23] ) | (~new_n507_ & (~new_n495_ | ~\a[23] ) & (new_n495_ | \a[23] )))) | ((new_n508_ ^ ~\a[23] ) & (~new_n495_ | ~\a[23] ) & (new_n507_ | (new_n495_ & \a[23] ) | (~new_n495_ & ~\a[23] )))) & (\a[20]  | ((~new_n508_ ^ ~\a[23] ) ^ ((new_n495_ & \a[23] ) | (~new_n507_ & (~new_n495_ | ~\a[23] ) & (new_n495_ | \a[23] )))))));
  assign new_n563_ = ((\a[20]  & (new_n507_ | (new_n495_ & \a[23] ) | (~new_n495_ & ~\a[23] )) & (~new_n507_ | (new_n495_ ^ \a[23] ))) | (~new_n69_ & (~\a[20]  | (~new_n507_ & (~new_n495_ | ~\a[23] ) & (new_n495_ | \a[23] )) | (new_n507_ & (~new_n495_ ^ \a[23] ))) & (\a[20]  | (~new_n507_ ^ (new_n495_ ^ \a[23] ))))) ^ (\a[20]  ^ ((new_n508_ ^ \a[23] ) ^ ((new_n495_ & \a[23] ) | (~new_n507_ & (~new_n495_ | ~\a[23] ) & (new_n495_ | \a[23] )))));
  assign new_n564_ = (~\a[17]  | (new_n69_ & ~new_n565_) | (~new_n69_ & new_n565_)) & ((\a[17]  & (~new_n69_ | new_n565_) & (new_n69_ | ~new_n565_)) | (~\a[17]  & (~new_n69_ ^ ~new_n565_)) | ((~new_n566_ | ~\a[17] ) & ((new_n566_ & \a[17] ) | (~new_n566_ & ~\a[17] ) | ((~new_n567_ | ~\a[17] ) & ((new_n567_ & \a[17] ) | (~new_n567_ & ~\a[17] ) | (~new_n568_ & (new_n569_ | ~new_n639_)))))));
  assign new_n565_ = \a[20]  ^ (~new_n507_ ^ (~new_n495_ ^ ~\a[23] ));
  assign new_n566_ = ((\a[20]  & ((new_n70_ & \a[23] ) | (~new_n70_ & ~\a[23] ) | ((~new_n361_ | ~\a[23] ) & ((new_n361_ & \a[23] ) | (~new_n361_ & ~\a[23] ) | ((~new_n362_ | ~\a[23] ) & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )))))) & ((new_n70_ ^ \a[23] ) | (new_n361_ & \a[23] ) | ((~new_n361_ | ~\a[23] ) & (new_n361_ | \a[23] ) & ((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )))))) | (((\a[20]  & ((new_n361_ & \a[23] ) | (~new_n361_ & ~\a[23] ) | ((~new_n362_ | ~\a[23] ) & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )))) & ((new_n361_ ^ \a[23] ) | (new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )))) | ((~\a[20]  | ((~new_n361_ | ~\a[23] ) & (new_n361_ | \a[23] ) & ((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )))) | ((~new_n361_ ^ \a[23] ) & (~new_n362_ | ~\a[23] ) & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )))) & (\a[20]  | ((new_n361_ ^ \a[23] ) ^ ((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] ))))) & ((\a[20]  & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )) & (~new_n363_ | (new_n362_ ^ \a[23] ))) | (~new_n429_ & (~\a[20]  | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )) | (new_n363_ & (~new_n362_ ^ \a[23] ))) & (\a[20]  | (~new_n363_ ^ (new_n362_ ^ \a[23] ))))))) & (~\a[20]  | ((~new_n70_ | ~\a[23] ) & (new_n70_ | \a[23] ) & ((new_n361_ & \a[23] ) | ((~new_n361_ | ~\a[23] ) & (new_n361_ | \a[23] ) & ((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )))))) | ((~new_n70_ ^ \a[23] ) & (~new_n361_ | ~\a[23] ) & ((new_n361_ & \a[23] ) | (~new_n361_ & ~\a[23] ) | ((~new_n362_ | ~\a[23] ) & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )))))) & (\a[20]  | ((new_n70_ ^ \a[23] ) ^ ((new_n361_ & \a[23] ) | ((~new_n361_ | ~\a[23] ) & (new_n361_ | \a[23] ) & ((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] ))))))))) ^ (new_n344_ ^ \a[20] );
  assign new_n567_ = ((\a[20]  & ((new_n361_ & \a[23] ) | (~new_n361_ & ~\a[23] ) | ((~new_n362_ | ~\a[23] ) & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )))) & ((new_n361_ ^ \a[23] ) | (new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )))) | (((\a[20]  & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )) & (~new_n363_ | (new_n362_ ^ \a[23] ))) | (~new_n429_ & (~\a[20]  | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )) | (new_n363_ & (~new_n362_ ^ \a[23] ))) & (\a[20]  | (~new_n363_ ^ (new_n362_ ^ \a[23] ))))) & (~\a[20]  | ((~new_n361_ | ~\a[23] ) & (new_n361_ | \a[23] ) & ((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )))) | ((~new_n361_ ^ \a[23] ) & (~new_n362_ | ~\a[23] ) & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )))) & (\a[20]  | ((new_n361_ ^ \a[23] ) ^ ((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] ))))))) ^ (\a[20]  ^ ((~new_n70_ ^ ~\a[23] ) ^ ((new_n361_ & \a[23] ) | ((~new_n361_ | ~\a[23] ) & (new_n361_ | \a[23] ) & ((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )))))));
  assign new_n568_ = \a[17]  & (((~\a[20]  | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )) | (new_n363_ & (~new_n362_ ^ \a[23] ))) & (new_n429_ | (\a[20]  & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )) & (~new_n363_ | (new_n362_ ^ \a[23] ))) | (~\a[20]  & (new_n363_ ^ (new_n362_ ^ \a[23] ))))) | (\a[20]  & (((~new_n362_ | ~\a[23] ) & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] ))) | (new_n361_ & \a[23] ) | (~new_n361_ & ~\a[23] )) & ((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )) | (new_n361_ ^ \a[23] ))) | (~\a[20]  & (((~new_n362_ | ~\a[23] ) & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] ))) ^ (new_n361_ ^ \a[23] )))) & ((\a[20]  & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )) & (~new_n363_ | (new_n362_ ^ \a[23] ))) | (~new_n429_ & (~\a[20]  | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )) | (new_n363_ & (~new_n362_ ^ \a[23] ))) & (\a[20]  | (~new_n363_ ^ (new_n362_ ^ \a[23] )))) | (\a[20]  ^ (((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] ))) ^ (new_n361_ ^ \a[23] ))));
  assign new_n569_ = (~\a[17]  | (new_n429_ & ~new_n570_) | (~new_n429_ & new_n570_)) & (((~new_n571_ | ~\a[17] ) & ((new_n571_ & \a[17] ) | (~new_n571_ & ~\a[17] ) | ((~new_n572_ | ~\a[17] ) & (((~new_n573_ | ~\a[17] ) & (new_n575_ | (~new_n573_ & ~\a[17] ) | (new_n573_ & \a[17] ))) | (new_n572_ & \a[17] ) | (~new_n572_ & ~\a[17] ))))) | (\a[17]  & (~new_n429_ | new_n570_) & (new_n429_ | ~new_n570_)) | (~\a[17]  & (~new_n429_ ^ ~new_n570_)));
  assign new_n570_ = \a[20]  ^ (~new_n363_ ^ (~new_n362_ ^ ~\a[23] ));
  assign new_n571_ = (~new_n430_ ^ ~\a[20] ) ^ ((\a[20]  & ((new_n365_ & \a[23] ) | (~new_n365_ & ~\a[23] ) | ((~new_n367_ | ~\a[23] ) & ((new_n367_ & \a[23] ) | (~new_n367_ & ~\a[23] ) | ((~new_n368_ | ~\a[23] ) & (new_n370_ | (new_n368_ & \a[23] ) | (~new_n368_ & ~\a[23] )))))) & ((new_n365_ ^ \a[23] ) | (new_n367_ & \a[23] ) | ((~new_n367_ | ~\a[23] ) & (new_n367_ | \a[23] ) & ((new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] )))))) | (((\a[20]  & ((new_n367_ & \a[23] ) | (~new_n367_ & ~\a[23] ) | ((~new_n368_ | ~\a[23] ) & (new_n370_ | (new_n368_ & \a[23] ) | (~new_n368_ & ~\a[23] )))) & ((new_n367_ ^ \a[23] ) | (new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] )))) | (~new_n431_ & (~\a[20]  | ((~new_n367_ | ~\a[23] ) & (new_n367_ | \a[23] ) & ((new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] )))) | ((~new_n367_ ^ \a[23] ) & (~new_n368_ | ~\a[23] ) & (new_n370_ | (new_n368_ & \a[23] ) | (~new_n368_ & ~\a[23] )))) & (\a[20]  | ((new_n367_ ^ \a[23] ) ^ ((new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] ))))))) & (~\a[20]  | ((~new_n365_ | ~\a[23] ) & (new_n365_ | \a[23] ) & ((new_n367_ & \a[23] ) | ((~new_n367_ | ~\a[23] ) & (new_n367_ | \a[23] ) & ((new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] )))))) | ((~new_n365_ ^ \a[23] ) & (~new_n367_ | ~\a[23] ) & ((new_n367_ & \a[23] ) | (~new_n367_ & ~\a[23] ) | ((~new_n368_ | ~\a[23] ) & (new_n370_ | (new_n368_ & \a[23] ) | (~new_n368_ & ~\a[23] )))))) & (\a[20]  | ((new_n365_ ^ \a[23] ) ^ ((new_n367_ & \a[23] ) | ((~new_n367_ | ~\a[23] ) & (new_n367_ | \a[23] ) & ((new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] )))))))));
  assign new_n572_ = ((\a[20]  & ((new_n367_ & \a[23] ) | (~new_n367_ & ~\a[23] ) | ((~new_n368_ | ~\a[23] ) & (new_n370_ | (new_n368_ & \a[23] ) | (~new_n368_ & ~\a[23] )))) & ((new_n367_ ^ \a[23] ) | (new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] )))) | (~new_n431_ & (~\a[20]  | ((~new_n367_ | ~\a[23] ) & (new_n367_ | \a[23] ) & ((new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] )))) | ((~new_n367_ ^ \a[23] ) & (~new_n368_ | ~\a[23] ) & (new_n370_ | (new_n368_ & \a[23] ) | (~new_n368_ & ~\a[23] )))) & (\a[20]  | ((new_n367_ ^ \a[23] ) ^ ((new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] ))))))) ^ (\a[20]  ^ ((new_n365_ ^ \a[23] ) ^ ((new_n367_ & \a[23] ) | ((~new_n367_ | ~\a[23] ) & (new_n367_ | \a[23] ) & ((new_n368_ & \a[23] ) | (~new_n370_ & (~new_n368_ | ~\a[23] ) & (new_n368_ | \a[23] )))))));
  assign new_n573_ = new_n431_ ^ ~new_n574_;
  assign new_n574_ = \a[20]  ^ ((new_n367_ ^ \a[23] ) ^ ((new_n368_ & \a[23] ) | (~new_n370_ & (new_n368_ | \a[23] ) & (~new_n368_ | ~\a[23] ))));
  assign new_n575_ = (~new_n576_ | ~\a[17] ) & ((~new_n576_ & ~\a[17] ) | (new_n576_ & \a[17] ) | ((~\a[17]  | ((~new_n433_ | ~\a[20] ) & (new_n433_ | \a[20] ) & ((new_n434_ & \a[20] ) | ((~new_n434_ | ~\a[20] ) & (new_n434_ | \a[20] ) & ((new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] )))))) | ((~new_n433_ ^ \a[20] ) & (~new_n434_ | ~\a[20] ) & ((new_n434_ & \a[20] ) | (~new_n434_ & ~\a[20] ) | ((~new_n435_ | ~\a[20] ) & (new_n436_ | (new_n435_ & \a[20] ) | (~new_n435_ & ~\a[20] )))))) & (((~\a[17]  | ((~new_n434_ | ~\a[20] ) & (new_n434_ | \a[20] ) & ((new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] )))) | ((~new_n434_ ^ \a[20] ) & (~new_n435_ | ~\a[20] ) & (new_n436_ | (new_n435_ & \a[20] ) | (~new_n435_ & ~\a[20] )))) & (new_n577_ | (\a[17]  & ((new_n434_ & \a[20] ) | (~new_n434_ & ~\a[20] ) | ((~new_n435_ | ~\a[20] ) & (new_n436_ | (new_n435_ & \a[20] ) | (~new_n435_ & ~\a[20] )))) & ((new_n434_ ^ \a[20] ) | (new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] )))) | (~\a[17]  & ((~new_n434_ ^ \a[20] ) ^ ((new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] ))))))) | (\a[17]  & ((new_n433_ & \a[20] ) | (~new_n433_ & ~\a[20] ) | ((~new_n434_ | ~\a[20] ) & ((new_n434_ & \a[20] ) | (~new_n434_ & ~\a[20] ) | ((~new_n435_ | ~\a[20] ) & (new_n436_ | (new_n435_ & \a[20] ) | (~new_n435_ & ~\a[20] )))))) & ((new_n433_ ^ \a[20] ) | (new_n434_ & \a[20] ) | ((~new_n434_ | ~\a[20] ) & (new_n434_ | \a[20] ) & ((new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] )))))) | (~\a[17]  & ((~new_n433_ ^ \a[20] ) ^ ((new_n434_ & \a[20] ) | ((~new_n434_ | ~\a[20] ) & (new_n434_ | \a[20] ) & ((new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] ))))))))));
  assign new_n576_ = ((new_n433_ & \a[20] ) | ((~new_n433_ | ~\a[20] ) & (new_n433_ | \a[20] ) & ((new_n434_ & \a[20] ) | (((new_n435_ & \a[20] ) | (~new_n436_ & (new_n435_ | \a[20] ) & (~new_n435_ | ~\a[20] ))) & (~new_n434_ | ~\a[20] ) & (new_n434_ | \a[20] ))))) ^ (\a[20]  ^ (new_n370_ ^ ~new_n432_));
  assign new_n577_ = (~\a[17]  | ((~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] ) & ((new_n437_ & \a[20] ) | (~new_n578_ & (~new_n437_ | ~\a[20] ) & (new_n437_ | \a[20] )))) | ((~new_n435_ ^ \a[20] ) & (~new_n437_ | ~\a[20] ) & (new_n578_ | (new_n437_ & \a[20] ) | (~new_n437_ & ~\a[20] )))) & (((~\a[17]  | (~new_n578_ & (~new_n437_ | ~\a[20] ) & (new_n437_ | \a[20] )) | (new_n578_ & (~new_n437_ ^ \a[20] ))) & (((~new_n579_ | ~\a[17] ) & ((new_n579_ & \a[17] ) | (~new_n579_ & ~\a[17] ) | ((~new_n580_ | ~\a[17] ) & (new_n581_ | (new_n580_ & \a[17] ) | (~new_n580_ & ~\a[17] ))))) | (\a[17]  & (new_n578_ | (new_n437_ & \a[20] ) | (~new_n437_ & ~\a[20] )) & (~new_n578_ | (new_n437_ ^ \a[20] ))) | (~\a[17]  & (new_n578_ ^ (new_n437_ ^ \a[20] ))))) | (\a[17]  & ((new_n435_ & \a[20] ) | (~new_n435_ & ~\a[20] ) | ((~new_n437_ | ~\a[20] ) & (new_n578_ | (new_n437_ & \a[20] ) | (~new_n437_ & ~\a[20] )))) & ((new_n435_ ^ \a[20] ) | (new_n437_ & \a[20] ) | (~new_n578_ & (~new_n437_ | ~\a[20] ) & (new_n437_ | \a[20] )))) | (~\a[17]  & ((~new_n435_ ^ \a[20] ) ^ ((new_n437_ & \a[20] ) | (~new_n578_ & (~new_n437_ | ~\a[20] ) & (new_n437_ | \a[20] ))))));
  assign new_n578_ = ~new_n438_ & (new_n438_ | new_n492_ | ((new_n493_ | (~new_n382_ & new_n423_) | (new_n382_ & ~new_n423_)) & (new_n440_ | (~new_n493_ & (new_n382_ | ~new_n423_) & (~new_n382_ | new_n423_)) | (new_n493_ & (new_n382_ ^ new_n423_)))));
  assign new_n579_ = (~new_n438_ & ~new_n492_) ^ ((~new_n493_ & (new_n382_ | ~new_n423_) & (~new_n382_ | new_n423_)) | (~new_n440_ & (new_n493_ | (~new_n382_ & new_n423_) | (new_n382_ & ~new_n423_)) & (~new_n493_ | (~new_n382_ ^ new_n423_))));
  assign new_n580_ = ~new_n440_ ^ (~new_n493_ ^ (~new_n382_ ^ new_n423_));
  assign new_n581_ = (~new_n582_ | ~\a[17] ) & ((new_n582_ & \a[17] ) | (~new_n582_ & ~\a[17] ) | (~new_n583_ & (new_n637_ | ((new_n638_ | (~new_n448_ & new_n489_) | (new_n448_ & ~new_n489_)) & (new_n585_ | (~new_n638_ & (new_n448_ | ~new_n489_) & (~new_n448_ | new_n489_)) | (new_n638_ & (new_n448_ ^ new_n489_)))))));
  assign new_n582_ = (new_n441_ ^ ~new_n491_) ^ (new_n443_ | (new_n490_ & (new_n445_ | (~new_n448_ & new_n489_))));
  assign new_n583_ = ~new_n584_ & (~new_n490_ | (~new_n445_ & (new_n448_ | ~new_n489_))) & (new_n490_ | new_n445_ | (~new_n448_ & new_n489_));
  assign new_n584_ = \a[17]  ^ (~\b[19]  | (((\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (new_n201_ | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ))));
  assign new_n585_ = (~new_n586_ | new_n636_) & ((new_n586_ & ~new_n636_) | (~new_n586_ & new_n636_) | (~new_n588_ & (~new_n635_ | (~new_n590_ & (new_n593_ | ~new_n634_)))));
  assign new_n586_ = new_n587_ ^ (new_n450_ | (((~new_n488_ & (new_n394_ | ~new_n417_) & (~new_n394_ | new_n417_)) | (~new_n452_ & (new_n488_ | (~new_n394_ & new_n417_) | (new_n394_ & ~new_n417_)) & (~new_n488_ | (~new_n394_ ^ new_n417_)))) & ~new_n450_ & ~new_n486_));
  assign new_n587_ = ~new_n487_ ^ ((new_n389_ | (new_n418_ & (new_n391_ | (~new_n394_ & new_n417_)))) ^ (new_n387_ ^ ~new_n419_));
  assign new_n588_ = ~new_n589_ & (new_n450_ | new_n486_ | ((new_n488_ | (~new_n394_ & new_n417_) | (new_n394_ & ~new_n417_)) & (new_n452_ | (~new_n488_ & (new_n394_ | ~new_n417_) & (~new_n394_ | new_n417_)) | (new_n488_ & (new_n394_ ^ new_n417_))))) & ((~new_n450_ & ~new_n486_) | (~new_n488_ & (new_n394_ | ~new_n417_) & (~new_n394_ | new_n417_)) | (~new_n452_ & (new_n488_ | (~new_n394_ & new_n417_) | (new_n394_ & ~new_n417_)) & (~new_n488_ | (~new_n394_ ^ new_n417_))));
  assign new_n589_ = \a[17]  ^ ((~\b[16]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[17]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[18]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  ^ \a[17] )) & (~new_n199_ | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )));
  assign new_n590_ = ~new_n592_ & (~new_n452_ | new_n591_) & (new_n452_ | ~new_n591_);
  assign new_n591_ = ~new_n488_ ^ (new_n394_ ^ ~new_n417_);
  assign new_n592_ = \a[17]  ^ ((~\b[15]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[16]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[17]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  ^ \a[17] )) & (~new_n144_ | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )));
  assign new_n593_ = (~new_n594_ | new_n632_) & ((new_n594_ & ~new_n632_) | (~new_n594_ & new_n632_) | (~new_n595_ & (new_n595_ | new_n631_ | ((new_n633_ | (~new_n460_ & new_n483_) | (new_n460_ & ~new_n483_)) & (new_n597_ | (~new_n633_ & (new_n460_ | ~new_n483_) & (~new_n460_ | new_n483_)) | (new_n633_ & (new_n460_ ^ new_n483_)))))));
  assign new_n594_ = (new_n453_ ^ ~new_n485_) ^ (new_n455_ | (new_n484_ & (new_n457_ | (~new_n460_ & new_n483_))));
  assign new_n595_ = ~new_n596_ & (~new_n484_ | (~new_n457_ & (new_n460_ | ~new_n483_))) & (new_n484_ | new_n457_ | (~new_n460_ & new_n483_));
  assign new_n596_ = \a[17]  ^ ((((~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] ) & ((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )))) | ((~\b[14]  ^ \b[15] ) & (~\b[13]  | ~\b[14] ) & (new_n142_ | (\b[13]  & \b[14] ) | (~\b[13]  & ~\b[14] ))) | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )) & (~\b[13]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[14]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[15]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  ^ \a[17] )));
  assign new_n597_ = (~new_n598_ | new_n630_) & ((new_n598_ & ~new_n630_) | (~new_n598_ & new_n630_) | (~new_n600_ & (~new_n629_ | (~new_n602_ & (new_n605_ | ~new_n628_)))));
  assign new_n598_ = new_n599_ ^ (new_n463_ | (new_n479_ & ((~new_n482_ & (new_n405_ | (~new_n404_ & new_n412_) | (new_n404_ & ~new_n412_)) & (~new_n405_ | (~new_n404_ ^ new_n412_))) | (~new_n465_ & (new_n482_ | (~new_n405_ & (new_n404_ | ~new_n412_) & (~new_n404_ | new_n412_)) | (new_n405_ & (new_n404_ ^ new_n412_))) & (~new_n482_ | (~new_n405_ ^ (~new_n404_ ^ new_n412_)))))));
  assign new_n599_ = ~new_n480_ ^ ((new_n400_ ^ ~new_n401_) ^ ((new_n402_ & ~new_n403_) | ((~new_n402_ | new_n403_) & (new_n402_ | ~new_n403_) & ((~new_n404_ & new_n412_) | (~new_n405_ & (new_n404_ | ~new_n412_) & (~new_n404_ | new_n412_))))));
  assign new_n600_ = ~new_n601_ & (~new_n479_ | ((new_n482_ | (~new_n405_ & (new_n404_ | ~new_n412_) & (~new_n404_ | new_n412_)) | (new_n405_ & (new_n404_ ^ new_n412_))) & (new_n465_ | (~new_n482_ & (new_n405_ | (~new_n404_ & new_n412_) | (new_n404_ & ~new_n412_)) & (~new_n405_ | (~new_n404_ ^ new_n412_))) | (new_n482_ & (new_n405_ ^ (~new_n404_ ^ new_n412_)))))) & (new_n479_ | (~new_n482_ & (new_n405_ | (~new_n404_ & new_n412_) | (new_n404_ & ~new_n412_)) & (~new_n405_ | (~new_n404_ ^ new_n412_))) | (~new_n465_ & (new_n482_ | (~new_n405_ & (new_n404_ | ~new_n412_) & (~new_n404_ | new_n412_)) | (new_n405_ & (new_n404_ ^ new_n412_))) & (~new_n482_ | (~new_n405_ ^ (~new_n404_ ^ new_n412_)))));
  assign new_n601_ = \a[17]  ^ ((~\b[10]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[11]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[12]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  ^ \a[17] )) & (~new_n107_ | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )));
  assign new_n602_ = ~new_n604_ & (~new_n465_ | new_n603_) & (new_n465_ | ~new_n603_);
  assign new_n603_ = ~new_n482_ ^ (~new_n405_ ^ (~new_n404_ ^ new_n412_));
  assign new_n604_ = \a[17]  ^ ((~\b[9]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[10]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[11]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  ^ \a[17] )) & (~new_n135_ | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )));
  assign new_n605_ = (~new_n607_ | new_n625_) & ((~new_n608_ & (~new_n624_ | ((new_n627_ | (new_n606_ & ~new_n471_) | (~new_n606_ & new_n471_)) & (new_n610_ | (~new_n627_ & (~new_n606_ | new_n471_) & (new_n606_ | ~new_n471_)) | (new_n627_ & (~new_n606_ ^ ~new_n471_)))))) | (new_n607_ & ~new_n625_) | (~new_n607_ & new_n625_));
  assign new_n606_ = new_n470_ ^ ~new_n478_;
  assign new_n607_ = (new_n466_ ^ ~new_n467_) ^ ((new_n468_ & ~new_n469_) | (((~new_n470_ & new_n478_) | (~new_n471_ & (new_n470_ | ~new_n478_) & (~new_n470_ | new_n478_))) & (~new_n468_ | new_n469_) & (new_n468_ | ~new_n469_)));
  assign new_n608_ = ~new_n609_ & ((new_n468_ & ~new_n469_) | (~new_n468_ & new_n469_) | ((new_n470_ | ~new_n478_) & (new_n471_ | (~new_n470_ & new_n478_) | (new_n470_ & ~new_n478_)))) & ((new_n468_ ^ ~new_n469_) | (~new_n470_ & new_n478_) | (~new_n471_ & (new_n470_ | ~new_n478_) & (~new_n470_ | new_n478_)));
  assign new_n609_ = \a[17]  ^ ((((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))) | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )) & (~\b[7]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[8]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[9]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  ^ \a[17] )));
  assign new_n610_ = (new_n611_ | ~new_n612_) & ((new_n611_ & ~new_n612_) | (~new_n611_ & new_n612_) | ((~new_n613_ | new_n614_) & (((new_n615_ | ~new_n623_) & (new_n616_ | (~new_n615_ & new_n623_) | (new_n615_ & ~new_n623_))) | (new_n613_ & ~new_n614_) | (~new_n613_ & new_n614_))));
  assign new_n611_ = \a[17]  ^ ((~\b[5]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[6]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[7]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  ^ \a[17] )) & (~new_n88_ | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )));
  assign new_n612_ = (new_n475_ | (~new_n476_ & new_n477_)) ^ (new_n474_ ^ (~\a[20]  ^ (new_n473_ & (~new_n98_ | ~new_n472_))));
  assign new_n613_ = new_n476_ ^ ~new_n477_;
  assign new_n614_ = \a[17]  ^ ((~\b[4]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[5]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[6]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  ^ \a[17] )) & (~new_n91_ | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )));
  assign new_n615_ = \a[17]  ^ ((~\b[3]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[4]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[5]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  ^ \a[17] )) & (~new_n94_ | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )));
  assign new_n616_ = (~new_n619_ | (\a[17]  ^ (new_n618_ & (~new_n98_ | ~new_n617_)))) & ((~new_n620_ & (new_n621_ | ~new_n622_)) | (new_n619_ & (~\a[17]  ^ (new_n618_ & (~new_n98_ | ~new_n617_)))) | (~new_n619_ & (~\a[17]  | ~new_n618_ | (new_n98_ & new_n617_)) & (\a[17]  | (new_n618_ & (~new_n98_ | ~new_n617_)))));
  assign new_n617_ = (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ) & (~\a[16]  | ~\a[17] ) & (\a[16]  | \a[17] );
  assign new_n618_ = (~\b[2]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[3]  | (~\a[14]  ^ ~\a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[4]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  ^ \a[17] ));
  assign new_n619_ = ((\b[0]  & (\a[17]  ^ ~\a[18] ) & (~\a[18]  | ~\a[19] ) & (\a[18]  | \a[19] )) | (\b[1]  & (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ) & (~\a[19]  ^ \a[20] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ) & (~\a[19]  | ~\a[20] ) & (\a[19]  | \a[20] ))) ^ (\a[20]  & \b[0]  & (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] ));
  assign new_n620_ = \b[0]  & (~\a[17]  | ~\a[18] ) & (\a[17]  | \a[18] ) & (~\b[0]  | (~\a[14]  ^ ~\a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[1]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  ^ \a[17] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )) & \a[17]  & (~\b[0]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[0]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[1]  | (~\a[14]  ^ ~\a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[2]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  ^ \a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )));
  assign new_n621_ = \a[17]  ^ (((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[2]  | (~\a[14]  ^ ~\a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[3]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  ^ \a[17] )));
  assign new_n622_ = (\b[0]  & (~\a[17]  | ~\a[18] ) & (\a[17]  | \a[18] )) ^ ((~\b[0]  | (~\a[14]  ^ ~\a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[1]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  ^ \a[17] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )) & \a[17]  & (~\b[0]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[0]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[1]  | (~\a[14]  ^ ~\a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[2]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  ^ \a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n623_ = ((~\b[0]  | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (~\a[17]  ^ ~\a[18] ) | (\a[18]  ^ \a[19] )) & (~\b[1]  | (~\a[17]  ^ ~\a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[2]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  ^ \a[20] )) & ((~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))) ^ (~\a[20]  | ((~\b[0]  | (~\a[17]  ^ ~\a[18] ) | (\a[18]  & \a[19] ) | (~\a[18]  & ~\a[19] )) & (~\b[1]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  ^ \a[20] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ) | (\a[19]  & \a[20] ) | (~\a[19]  & ~\a[20] )) & \a[20]  & (~\b[0]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ))));
  assign new_n624_ = ~new_n609_ ^ ((new_n468_ ^ ~new_n469_) ^ ((~new_n470_ & new_n478_) | (~new_n471_ & (new_n470_ | ~new_n478_) & (~new_n470_ | new_n478_))));
  assign new_n625_ = \a[17]  ^ (new_n626_ & (~new_n617_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n626_ = (~\b[8]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[9]  | (~\a[14]  ^ ~\a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[10]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  ^ \a[17] ));
  assign new_n627_ = \a[17]  ^ ((~\b[6]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[7]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[8]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  ^ \a[17] )) & ((\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n79_ & (~\b[7]  ^ \b[8] ))));
  assign new_n628_ = ~new_n604_ ^ (new_n465_ ^ ~new_n603_);
  assign new_n629_ = ~new_n601_ ^ (new_n479_ ^ ((~new_n482_ & (new_n405_ | (~new_n404_ & new_n412_) | (new_n404_ & ~new_n412_)) & (~new_n405_ | (~new_n404_ ^ new_n412_))) | (~new_n465_ & (new_n482_ | (~new_n405_ & (new_n404_ | ~new_n412_) & (~new_n404_ | new_n412_)) | (new_n405_ & (new_n404_ ^ new_n412_))) & (~new_n482_ | (~new_n405_ ^ (~new_n404_ ^ new_n412_))))));
  assign new_n630_ = \a[17]  ^ ((~\b[11]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[12]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[13]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  ^ \a[17] )) & (~new_n133_ | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )));
  assign new_n631_ = new_n596_ & (~new_n484_ ^ (new_n457_ | (~new_n460_ & new_n483_)));
  assign new_n632_ = \a[17]  ^ ((~\b[14]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[15]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[16]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  ^ \a[17] )) & (~new_n186_ | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )));
  assign new_n633_ = \a[17]  ^ ((~\b[12]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[13]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[14]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  ^ \a[17] )) & ((\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n142_ & (~\b[13]  ^ \b[14] ))));
  assign new_n634_ = ~new_n592_ ^ (new_n452_ ^ ~new_n591_);
  assign new_n635_ = ~new_n589_ ^ ((~new_n450_ & ~new_n486_) ^ ((~new_n488_ & (new_n394_ | ~new_n417_) & (~new_n394_ | new_n417_)) | (~new_n452_ & (new_n488_ | (~new_n394_ & new_n417_) | (new_n394_ & ~new_n417_)) & (~new_n488_ | (~new_n394_ ^ new_n417_)))));
  assign new_n636_ = \a[17]  ^ ((~\b[17]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[18]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[19]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  ^ \a[17] )) & (~new_n253_ | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )));
  assign new_n637_ = new_n584_ & (~new_n490_ ^ (new_n445_ | (~new_n448_ & new_n489_)));
  assign new_n638_ = \a[17]  ^ (((\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~new_n201_ ^ ~\b[19] )) & (~\b[18]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\a[14]  ^ \a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[19]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )));
  assign new_n639_ = \a[17]  ^ (((\a[20]  & (new_n363_ | (new_n362_ & \a[23] ) | (~new_n362_ & ~\a[23] )) & (~new_n363_ | (new_n362_ ^ \a[23] ))) | (~new_n429_ & (~\a[20]  | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] )) | (new_n363_ & (~new_n362_ ^ \a[23] ))) & (\a[20]  | (~new_n363_ ^ (new_n362_ ^ \a[23] ))))) ^ (\a[20]  ^ (((new_n362_ & \a[23] ) | (~new_n363_ & (~new_n362_ | ~\a[23] ) & (new_n362_ | \a[23] ))) ^ (new_n361_ ^ \a[23] ))));
  assign new_n640_ = (~new_n721_ | ~\a[8] ) & (((~\a[8]  | ((~new_n641_ | ~\a[11] ) & (new_n641_ | \a[11] ) & ((new_n723_ & \a[11] ) | ((~new_n723_ | ~\a[11] ) & (new_n723_ | \a[11] ) & ((new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] )))))) | ((~new_n641_ ^ \a[11] ) & (~new_n723_ | ~\a[11] ) & ((new_n723_ & \a[11] ) | (~new_n723_ & ~\a[11] ) | ((~new_n724_ | ~\a[11] ) & (new_n725_ | (new_n724_ & \a[11] ) | (~new_n724_ & ~\a[11] )))))) & (((~\a[8]  | ((~new_n723_ | ~\a[11] ) & (new_n723_ | \a[11] ) & ((new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] )))) | ((~new_n723_ ^ \a[11] ) & (~new_n724_ | ~\a[11] ) & (new_n725_ | (new_n724_ & \a[11] ) | (~new_n724_ & ~\a[11] )))) & ((\a[8]  & ((new_n723_ & \a[11] ) | (~new_n723_ & ~\a[11] ) | ((~new_n724_ | ~\a[11] ) & (new_n725_ | (new_n724_ & \a[11] ) | (~new_n724_ & ~\a[11] )))) & ((new_n723_ ^ \a[11] ) | (new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] )))) | (~\a[8]  & ((~new_n723_ ^ \a[11] ) ^ ((new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] ))))) | ((~\a[8]  | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] )) | (new_n725_ & (~new_n724_ ^ \a[11] ))) & (new_n807_ | (\a[8]  & (new_n725_ | (new_n724_ & \a[11] ) | (~new_n724_ & ~\a[11] )) & (~new_n725_ | (new_n724_ ^ \a[11] ))) | (~\a[8]  & (new_n725_ ^ (new_n724_ ^ \a[11] ))))))) | (\a[8]  & ((new_n641_ & \a[11] ) | (~new_n641_ & ~\a[11] ) | ((~new_n723_ | ~\a[11] ) & ((new_n723_ & \a[11] ) | (~new_n723_ & ~\a[11] ) | ((~new_n724_ | ~\a[11] ) & (new_n725_ | (new_n724_ & \a[11] ) | (~new_n724_ & ~\a[11] )))))) & ((new_n641_ ^ \a[11] ) | (new_n723_ & \a[11] ) | ((~new_n723_ | ~\a[11] ) & (new_n723_ | \a[11] ) & ((new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] )))))) | (~\a[8]  & ((~new_n641_ ^ \a[11] ) ^ ((new_n723_ & \a[11] ) | ((~new_n723_ | ~\a[11] ) & (new_n723_ | \a[11] ) & ((new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] ))))))))) | (new_n721_ & \a[8] ) | (~new_n721_ & ~\a[8] ));
  assign new_n641_ = ~new_n643_ ^ (~new_n642_ ^ ~\a[14] );
  assign new_n642_ = ~new_n564_ ^ (~new_n563_ ^ ~\a[17] );
  assign new_n643_ = (~\a[14]  | (new_n645_ & ((new_n566_ & \a[17] ) | (~new_n644_ & (~new_n566_ | ~\a[17] ) & (new_n566_ | \a[17] )))) | (~new_n645_ & (~new_n566_ | ~\a[17] ) & (new_n644_ | (new_n566_ & \a[17] ) | (~new_n566_ & ~\a[17] )))) & (((~\a[14]  | (~new_n644_ & (~new_n566_ | ~\a[17] ) & (new_n566_ | \a[17] )) | (new_n644_ & (~new_n566_ ^ \a[17] ))) & (((~new_n646_ | ~\a[14] ) & ((new_n646_ & \a[14] ) | (~new_n646_ & ~\a[14] ) | ((~new_n647_ | ~\a[14] ) & (new_n648_ | (new_n647_ & \a[14] ) | (~new_n647_ & ~\a[14] ))))) | (\a[14]  & (new_n644_ | (new_n566_ & \a[17] ) | (~new_n566_ & ~\a[17] )) & (~new_n644_ | (new_n566_ ^ \a[17] ))) | (~\a[14]  & (new_n644_ ^ (new_n566_ ^ \a[17] ))))) | (\a[14]  & (~new_n645_ | ((~new_n566_ | ~\a[17] ) & (new_n644_ | (new_n566_ & \a[17] ) | (~new_n566_ & ~\a[17] )))) & (new_n645_ | (new_n566_ & \a[17] ) | (~new_n644_ & (~new_n566_ | ~\a[17] ) & (new_n566_ | \a[17] )))) | (~\a[14]  & (~new_n645_ ^ ((new_n566_ & \a[17] ) | (~new_n644_ & (~new_n566_ | ~\a[17] ) & (new_n566_ | \a[17] ))))));
  assign new_n644_ = (~new_n567_ | ~\a[17] ) & ((~new_n568_ & (new_n569_ | ~new_n639_)) | (new_n567_ & \a[17] ) | (~new_n567_ & ~\a[17] ));
  assign new_n645_ = \a[17]  ^ (new_n69_ ^ ~new_n565_);
  assign new_n646_ = (new_n568_ | (~new_n569_ & new_n639_)) ^ (new_n567_ ^ \a[17] );
  assign new_n647_ = new_n569_ ^ ~new_n639_;
  assign new_n648_ = (~new_n649_ | ~\a[14] ) & ((~new_n649_ & ~\a[14] ) | (new_n649_ & \a[14] ) | ((~\a[14]  | ((~new_n571_ | ~\a[17] ) & (new_n571_ | \a[17] ) & ((new_n572_ & \a[17] ) | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))))) | ((~new_n571_ ^ \a[17] ) & (~new_n572_ | ~\a[17] ) & ((new_n572_ & \a[17] ) | (~new_n572_ & ~\a[17] ) | ((~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))))) & ((\a[14]  & ((new_n571_ & \a[17] ) | (~new_n571_ & ~\a[17] ) | ((~new_n572_ | ~\a[17] ) & ((new_n572_ & \a[17] ) | (~new_n572_ & ~\a[17] ) | ((~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))))) & ((new_n571_ ^ \a[17] ) | (new_n572_ & \a[17] ) | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))))) | (~\a[14]  & ((~new_n571_ ^ \a[17] ) ^ ((new_n572_ & \a[17] ) | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] ))))))) | ((~\a[14]  | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))) | ((~new_n572_ ^ \a[17] ) & (~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))) & ((\a[14]  & ((new_n572_ & \a[17] ) | (~new_n572_ & ~\a[17] ) | ((~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))) & ((new_n572_ ^ \a[17] ) | (new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))) | (~\a[14]  & ((~new_n572_ ^ \a[17] ) ^ ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] ))))) | ((~\a[14]  | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )) | (new_n575_ & (~new_n573_ ^ \a[17] ))) & (new_n650_ | (\a[14]  & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )) & (~new_n575_ | (new_n573_ ^ \a[17] ))) | (~\a[14]  & (new_n575_ ^ (new_n573_ ^ \a[17] ))))))))));
  assign new_n649_ = ((new_n571_ & \a[17] ) | ((~new_n571_ | ~\a[17] ) & (new_n571_ | \a[17] ) & ((new_n572_ & \a[17] ) | (((new_n573_ & \a[17] ) | (~new_n575_ & (new_n573_ | \a[17] ) & (~new_n573_ | ~\a[17] ))) & (~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ))))) ^ (\a[17]  ^ (new_n429_ ^ ~new_n570_));
  assign new_n650_ = (~new_n651_ | ~\a[14] ) & ((new_n651_ & \a[14] ) | (~new_n651_ & ~\a[14] ) | ((~new_n652_ | ~\a[14] ) & ((new_n652_ & \a[14] ) | (~new_n652_ & ~\a[14] ) | (~new_n653_ & (new_n655_ | ~new_n720_)))));
  assign new_n651_ = (~new_n576_ ^ ~\a[17] ) ^ ((\a[17]  & ((new_n433_ & \a[20] ) | (~new_n433_ & ~\a[20] ) | ((~new_n434_ | ~\a[20] ) & ((new_n434_ & \a[20] ) | (~new_n434_ & ~\a[20] ) | ((~new_n435_ | ~\a[20] ) & (new_n436_ | (new_n435_ & \a[20] ) | (~new_n435_ & ~\a[20] )))))) & ((new_n433_ ^ \a[20] ) | (new_n434_ & \a[20] ) | ((~new_n434_ | ~\a[20] ) & (new_n434_ | \a[20] ) & ((new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] )))))) | (((\a[17]  & ((new_n434_ & \a[20] ) | (~new_n434_ & ~\a[20] ) | ((~new_n435_ | ~\a[20] ) & (new_n436_ | (new_n435_ & \a[20] ) | (~new_n435_ & ~\a[20] )))) & ((new_n434_ ^ \a[20] ) | (new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] )))) | (~new_n577_ & (~\a[17]  | ((~new_n434_ | ~\a[20] ) & (new_n434_ | \a[20] ) & ((new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] )))) | ((~new_n434_ ^ \a[20] ) & (~new_n435_ | ~\a[20] ) & (new_n436_ | (new_n435_ & \a[20] ) | (~new_n435_ & ~\a[20] )))) & (\a[17]  | ((new_n434_ ^ \a[20] ) ^ ((new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] ))))))) & (~\a[17]  | ((~new_n433_ | ~\a[20] ) & (new_n433_ | \a[20] ) & ((new_n434_ & \a[20] ) | ((~new_n434_ | ~\a[20] ) & (new_n434_ | \a[20] ) & ((new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] )))))) | ((~new_n433_ ^ \a[20] ) & (~new_n434_ | ~\a[20] ) & ((new_n434_ & \a[20] ) | (~new_n434_ & ~\a[20] ) | ((~new_n435_ | ~\a[20] ) & (new_n436_ | (new_n435_ & \a[20] ) | (~new_n435_ & ~\a[20] )))))) & (\a[17]  | ((new_n433_ ^ \a[20] ) ^ ((new_n434_ & \a[20] ) | ((~new_n434_ | ~\a[20] ) & (new_n434_ | \a[20] ) & ((new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] )))))))));
  assign new_n652_ = ((\a[17]  & ((new_n434_ & \a[20] ) | (~new_n434_ & ~\a[20] ) | ((~new_n435_ | ~\a[20] ) & (new_n436_ | (new_n435_ & \a[20] ) | (~new_n435_ & ~\a[20] )))) & ((new_n434_ ^ \a[20] ) | (new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] )))) | (~new_n577_ & (~\a[17]  | ((~new_n434_ | ~\a[20] ) & (new_n434_ | \a[20] ) & ((new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] )))) | ((~new_n434_ ^ \a[20] ) & (~new_n435_ | ~\a[20] ) & (new_n436_ | (new_n435_ & \a[20] ) | (~new_n435_ & ~\a[20] )))) & (\a[17]  | ((new_n434_ ^ \a[20] ) ^ ((new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] ))))))) ^ (\a[17]  ^ ((new_n433_ ^ \a[20] ) ^ ((new_n434_ & \a[20] ) | ((~new_n434_ | ~\a[20] ) & (new_n434_ | \a[20] ) & ((new_n435_ & \a[20] ) | (~new_n436_ & (~new_n435_ | ~\a[20] ) & (new_n435_ | \a[20] )))))));
  assign new_n653_ = \a[14]  & (~new_n577_ | new_n654_) & (new_n577_ | ~new_n654_);
  assign new_n654_ = \a[17]  ^ ((new_n434_ ^ \a[20] ) ^ ((new_n435_ & \a[20] ) | (~new_n436_ & (new_n435_ | \a[20] ) & (~new_n435_ | ~\a[20] ))));
  assign new_n655_ = (~new_n657_ | ~\a[14] ) & ((new_n657_ & \a[14] ) | (~new_n657_ & ~\a[14] ) | ((~\a[14]  | ((~new_n656_ | ~\a[17] ) & (new_n656_ | \a[17] ) & ((new_n579_ & \a[17] ) | ((~new_n579_ | ~\a[17] ) & (new_n579_ | \a[17] ) & ((new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] )))))) | ((~new_n656_ ^ \a[17] ) & (~new_n579_ | ~\a[17] ) & ((new_n579_ & \a[17] ) | (~new_n579_ & ~\a[17] ) | ((~new_n580_ | ~\a[17] ) & (new_n581_ | (new_n580_ & \a[17] ) | (~new_n580_ & ~\a[17] )))))) & ((\a[14]  & ((new_n656_ & \a[17] ) | (~new_n656_ & ~\a[17] ) | ((~new_n579_ | ~\a[17] ) & ((new_n579_ & \a[17] ) | (~new_n579_ & ~\a[17] ) | ((~new_n580_ | ~\a[17] ) & (new_n581_ | (new_n580_ & \a[17] ) | (~new_n580_ & ~\a[17] )))))) & ((new_n656_ ^ \a[17] ) | (new_n579_ & \a[17] ) | ((~new_n579_ | ~\a[17] ) & (new_n579_ | \a[17] ) & ((new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] )))))) | (~\a[14]  & ((~new_n656_ ^ \a[17] ) ^ ((new_n579_ & \a[17] ) | ((~new_n579_ | ~\a[17] ) & (new_n579_ | \a[17] ) & ((new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] ))))))) | ((~\a[14]  | ((~new_n579_ | ~\a[17] ) & (new_n579_ | \a[17] ) & ((new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] )))) | ((~new_n579_ ^ \a[17] ) & (~new_n580_ | ~\a[17] ) & (new_n581_ | (new_n580_ & \a[17] ) | (~new_n580_ & ~\a[17] )))) & (new_n658_ | (\a[14]  & ((new_n579_ & \a[17] ) | (~new_n579_ & ~\a[17] ) | ((~new_n580_ | ~\a[17] ) & (new_n581_ | (new_n580_ & \a[17] ) | (~new_n580_ & ~\a[17] )))) & ((new_n579_ ^ \a[17] ) | (new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] )))) | (~\a[14]  & ((~new_n579_ ^ \a[17] ) ^ ((new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] ))))))))));
  assign new_n656_ = ~new_n578_ ^ (new_n437_ ^ \a[20] );
  assign new_n657_ = ((\a[17]  & (new_n578_ | (new_n437_ & \a[20] ) | (~new_n437_ & ~\a[20] )) & (~new_n578_ | (new_n437_ ^ \a[20] ))) | (((new_n579_ & \a[17] ) | ((~new_n579_ | ~\a[17] ) & (new_n579_ | \a[17] ) & ((new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] ))))) & (~\a[17]  | (~new_n578_ & (~new_n437_ | ~\a[20] ) & (new_n437_ | \a[20] )) | (new_n578_ & (~new_n437_ ^ \a[20] ))) & (\a[17]  | (~new_n578_ ^ (new_n437_ ^ \a[20] ))))) ^ (\a[17]  ^ ((new_n435_ ^ \a[20] ) ^ ((new_n437_ & \a[20] ) | (~new_n578_ & (~new_n437_ | ~\a[20] ) & (new_n437_ | \a[20] )))));
  assign new_n658_ = (~\a[14]  | ((~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] ) & ((new_n582_ & \a[17] ) | (~new_n659_ & (~new_n582_ | ~\a[17] ) & (new_n582_ | \a[17] )))) | ((~new_n580_ ^ \a[17] ) & (~new_n582_ | ~\a[17] ) & (new_n659_ | (new_n582_ & \a[17] ) | (~new_n582_ & ~\a[17] )))) & ((\a[14]  & ((new_n580_ & \a[17] ) | (~new_n580_ & ~\a[17] ) | ((~new_n582_ | ~\a[17] ) & (new_n659_ | (new_n582_ & \a[17] ) | (~new_n582_ & ~\a[17] )))) & ((new_n580_ ^ \a[17] ) | (new_n582_ & \a[17] ) | (~new_n659_ & (~new_n582_ | ~\a[17] ) & (new_n582_ | \a[17] )))) | (~\a[14]  & ((~new_n580_ ^ \a[17] ) ^ ((new_n582_ & \a[17] ) | (~new_n659_ & (~new_n582_ | ~\a[17] ) & (new_n582_ | \a[17] ))))) | ((~\a[14]  | (~new_n659_ & (~new_n582_ | ~\a[17] ) & (new_n582_ | \a[17] )) | (new_n659_ & (~new_n582_ ^ \a[17] ))) & ((\a[14]  & (new_n659_ | (new_n582_ & \a[17] ) | (~new_n582_ & ~\a[17] )) & (~new_n659_ | (new_n582_ ^ \a[17] ))) | (~\a[14]  & (new_n659_ ^ (new_n582_ ^ \a[17] ))) | ((new_n660_ | ~\a[14] ) & ((~new_n660_ & \a[14] ) | (new_n660_ & ~\a[14] ) | ((~new_n661_ | ~\a[14] ) & (new_n662_ | (new_n661_ & \a[14] ) | (~new_n661_ & ~\a[14] ))))))));
  assign new_n659_ = ~new_n583_ & (new_n637_ | ((new_n638_ | (~new_n448_ & new_n489_) | (new_n448_ & ~new_n489_)) & (new_n585_ | (~new_n638_ & (new_n448_ | ~new_n489_) & (~new_n448_ | new_n489_)) | (new_n638_ & (new_n448_ ^ new_n489_)))));
  assign new_n660_ = (~new_n583_ & ~new_n637_) ^ ((new_n638_ | (~new_n448_ & new_n489_) | (new_n448_ & ~new_n489_)) & (new_n585_ | (~new_n638_ & (new_n448_ | ~new_n489_) & (~new_n448_ | new_n489_)) | (new_n638_ & (new_n448_ ^ new_n489_))));
  assign new_n661_ = ~new_n585_ ^ (~new_n638_ ^ (~new_n448_ ^ new_n489_));
  assign new_n662_ = (~new_n663_ | ~\a[14] ) & ((new_n663_ & \a[14] ) | (~new_n663_ & ~\a[14] ) | (~new_n664_ & (new_n718_ | ((new_n719_ | (~new_n593_ & new_n634_) | (new_n593_ & ~new_n634_)) & (new_n666_ | (~new_n719_ & (new_n593_ | ~new_n634_) & (~new_n593_ | new_n634_)) | (new_n719_ & (new_n593_ ^ new_n634_)))))));
  assign new_n663_ = (new_n586_ ^ ~new_n636_) ^ (new_n588_ | (new_n635_ & (new_n590_ | (~new_n593_ & new_n634_))));
  assign new_n664_ = ~new_n665_ & (~new_n635_ | (~new_n590_ & (new_n593_ | ~new_n634_))) & (new_n635_ | new_n590_ | (~new_n593_ & new_n634_));
  assign new_n665_ = \a[14]  ^ (~\b[19]  | (((\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (new_n201_ | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ))));
  assign new_n666_ = (~new_n667_ | new_n717_) & ((new_n667_ & ~new_n717_) | (~new_n667_ & new_n717_) | (~new_n669_ & (~new_n716_ | (~new_n671_ & (new_n674_ | ~new_n715_)))));
  assign new_n667_ = new_n668_ ^ (new_n595_ | (((~new_n633_ & (new_n460_ | ~new_n483_) & (~new_n460_ | new_n483_)) | (~new_n597_ & (new_n633_ | (~new_n460_ & new_n483_) | (new_n460_ & ~new_n483_)) & (~new_n633_ | (~new_n460_ ^ new_n483_)))) & ~new_n595_ & ~new_n631_));
  assign new_n668_ = ~new_n632_ ^ ((new_n455_ | (new_n484_ & (new_n457_ | (~new_n460_ & new_n483_)))) ^ (new_n453_ ^ ~new_n485_));
  assign new_n669_ = ~new_n670_ & (new_n595_ | new_n631_ | ((new_n633_ | (~new_n460_ & new_n483_) | (new_n460_ & ~new_n483_)) & (new_n597_ | (~new_n633_ & (new_n460_ | ~new_n483_) & (~new_n460_ | new_n483_)) | (new_n633_ & (new_n460_ ^ new_n483_))))) & ((~new_n595_ & ~new_n631_) | (~new_n633_ & (new_n460_ | ~new_n483_) & (~new_n460_ | new_n483_)) | (~new_n597_ & (new_n633_ | (~new_n460_ & new_n483_) | (new_n460_ & ~new_n483_)) & (~new_n633_ | (~new_n460_ ^ new_n483_))));
  assign new_n670_ = \a[14]  ^ ((~\b[16]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[17]  | (\a[11]  ^ \a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[18]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  ^ \a[14] )) & (~new_n199_ | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n671_ = ~new_n673_ & (~new_n597_ | new_n672_) & (new_n597_ | ~new_n672_);
  assign new_n672_ = ~new_n633_ ^ (new_n460_ ^ ~new_n483_);
  assign new_n673_ = \a[14]  ^ ((~\b[15]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[16]  | (\a[11]  ^ \a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[17]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  ^ \a[14] )) & (~new_n144_ | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n674_ = (~new_n675_ | new_n713_) & ((new_n675_ & ~new_n713_) | (~new_n675_ & new_n713_) | (~new_n676_ & (new_n676_ | new_n712_ | ((new_n714_ | (~new_n605_ & new_n628_) | (new_n605_ & ~new_n628_)) & (new_n678_ | (~new_n714_ & (new_n605_ | ~new_n628_) & (~new_n605_ | new_n628_)) | (new_n714_ & (new_n605_ ^ new_n628_)))))));
  assign new_n675_ = (new_n598_ ^ ~new_n630_) ^ (new_n600_ | (new_n629_ & (new_n602_ | (~new_n605_ & new_n628_))));
  assign new_n676_ = ~new_n677_ & (~new_n629_ | (~new_n602_ & (new_n605_ | ~new_n628_))) & (new_n629_ | new_n602_ | (~new_n605_ & new_n628_));
  assign new_n677_ = \a[14]  ^ ((((~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] ) & ((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )))) | ((~\b[14]  ^ \b[15] ) & (~\b[13]  | ~\b[14] ) & (new_n142_ | (\b[13]  & \b[14] ) | (~\b[13]  & ~\b[14] ))) | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & (~\b[13]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[14]  | (\a[11]  ^ \a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[15]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  ^ \a[14] )));
  assign new_n678_ = (~new_n679_ | new_n711_) & ((new_n679_ & ~new_n711_) | (~new_n679_ & new_n711_) | (~new_n681_ & (~new_n710_ | (~new_n683_ & (new_n686_ | ~new_n709_)))));
  assign new_n679_ = new_n680_ ^ (new_n608_ | (new_n624_ & ((~new_n627_ & (new_n471_ | (~new_n470_ & new_n478_) | (new_n470_ & ~new_n478_)) & (~new_n471_ | (~new_n470_ ^ new_n478_))) | (~new_n610_ & (new_n627_ | (~new_n471_ & (new_n470_ | ~new_n478_) & (~new_n470_ | new_n478_)) | (new_n471_ & (new_n470_ ^ new_n478_))) & (~new_n627_ | (~new_n471_ ^ (~new_n470_ ^ new_n478_)))))));
  assign new_n680_ = ~new_n625_ ^ ((new_n466_ ^ ~new_n467_) ^ ((new_n468_ & ~new_n469_) | ((~new_n468_ | new_n469_) & (new_n468_ | ~new_n469_) & ((~new_n470_ & new_n478_) | (~new_n471_ & (new_n470_ | ~new_n478_) & (~new_n470_ | new_n478_))))));
  assign new_n681_ = ~new_n682_ & (~new_n624_ | ((new_n627_ | (~new_n471_ & (new_n470_ | ~new_n478_) & (~new_n470_ | new_n478_)) | (new_n471_ & (new_n470_ ^ new_n478_))) & (new_n610_ | (~new_n627_ & (new_n471_ | (~new_n470_ & new_n478_) | (new_n470_ & ~new_n478_)) & (~new_n471_ | (~new_n470_ ^ new_n478_))) | (new_n627_ & (new_n471_ ^ (~new_n470_ ^ new_n478_)))))) & (new_n624_ | (~new_n627_ & (new_n471_ | (~new_n470_ & new_n478_) | (new_n470_ & ~new_n478_)) & (~new_n471_ | (~new_n470_ ^ new_n478_))) | (~new_n610_ & (new_n627_ | (~new_n471_ & (new_n470_ | ~new_n478_) & (~new_n470_ | new_n478_)) | (new_n471_ & (new_n470_ ^ new_n478_))) & (~new_n627_ | (~new_n471_ ^ (~new_n470_ ^ new_n478_)))));
  assign new_n682_ = \a[14]  ^ ((~\b[10]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[11]  | (\a[11]  ^ \a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[12]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  ^ \a[14] )) & (~new_n107_ | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n683_ = ~new_n685_ & (~new_n610_ | new_n684_) & (new_n610_ | ~new_n684_);
  assign new_n684_ = ~new_n627_ ^ (~new_n471_ ^ (~new_n470_ ^ new_n478_));
  assign new_n685_ = \a[14]  ^ ((~\b[9]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[10]  | (\a[11]  ^ \a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[11]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  ^ \a[14] )) & (~new_n135_ | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n686_ = (~new_n688_ | new_n706_) & ((~new_n689_ & (~new_n705_ | ((new_n708_ | (new_n687_ & ~new_n616_) | (~new_n687_ & new_n616_)) & (new_n691_ | (~new_n708_ & (~new_n687_ | new_n616_) & (new_n687_ | ~new_n616_)) | (new_n708_ & (~new_n687_ ^ ~new_n616_)))))) | (new_n688_ & ~new_n706_) | (~new_n688_ & new_n706_));
  assign new_n687_ = new_n615_ ^ ~new_n623_;
  assign new_n688_ = (new_n611_ ^ ~new_n612_) ^ ((new_n613_ & ~new_n614_) | (((~new_n615_ & new_n623_) | (~new_n616_ & (new_n615_ | ~new_n623_) & (~new_n615_ | new_n623_))) & (~new_n613_ | new_n614_) & (new_n613_ | ~new_n614_)));
  assign new_n689_ = ~new_n690_ & ((new_n613_ & ~new_n614_) | (~new_n613_ & new_n614_) | ((new_n615_ | ~new_n623_) & (new_n616_ | (~new_n615_ & new_n623_) | (new_n615_ & ~new_n623_)))) & ((new_n613_ ^ ~new_n614_) | (~new_n615_ & new_n623_) | (~new_n616_ & (new_n615_ | ~new_n623_) & (~new_n615_ | new_n623_)));
  assign new_n690_ = \a[14]  ^ ((((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))) | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & (~\b[7]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[8]  | (\a[11]  ^ \a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[9]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  ^ \a[14] )));
  assign new_n691_ = (new_n692_ | ~new_n693_) & ((new_n692_ & ~new_n693_) | (~new_n692_ & new_n693_) | ((~new_n694_ | new_n695_) & (((new_n696_ | ~new_n704_) & (new_n697_ | (~new_n696_ & new_n704_) | (new_n696_ & ~new_n704_))) | (new_n694_ & ~new_n695_) | (~new_n694_ & new_n695_))));
  assign new_n692_ = \a[14]  ^ ((~\b[5]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[6]  | (\a[11]  ^ \a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[7]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  ^ \a[14] )) & (~new_n88_ | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n693_ = (new_n620_ | (~new_n621_ & new_n622_)) ^ (new_n619_ ^ (~\a[17]  ^ (new_n618_ & (~new_n98_ | ~new_n617_))));
  assign new_n694_ = new_n621_ ^ ~new_n622_;
  assign new_n695_ = \a[14]  ^ ((~\b[4]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[5]  | (\a[11]  ^ \a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[6]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  ^ \a[14] )) & (~new_n91_ | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n696_ = \a[14]  ^ ((~\b[3]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[4]  | (\a[11]  ^ \a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[5]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  ^ \a[14] )) & (~new_n94_ | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n697_ = (~new_n700_ | (\a[14]  ^ (new_n699_ & (~new_n98_ | ~new_n698_)))) & ((~new_n701_ & (new_n702_ | ~new_n703_)) | (new_n700_ & (~\a[14]  ^ (new_n699_ & (~new_n98_ | ~new_n698_)))) | (~new_n700_ & (~\a[14]  | ~new_n699_ | (new_n98_ & new_n698_)) & (\a[14]  | (new_n699_ & (~new_n98_ | ~new_n698_)))));
  assign new_n698_ = (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ) & (~\a[13]  | ~\a[14] ) & (\a[13]  | \a[14] );
  assign new_n699_ = (~\b[2]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[3]  | (~\a[11]  ^ ~\a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[4]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  ^ \a[14] ));
  assign new_n700_ = ((\b[0]  & (\a[14]  ^ ~\a[15] ) & (~\a[15]  | ~\a[16] ) & (\a[15]  | \a[16] )) | (\b[1]  & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ) & (~\a[16]  ^ \a[17] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ) & (~\a[16]  | ~\a[17] ) & (\a[16]  | \a[17] ))) ^ (\a[17]  & \b[0]  & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ));
  assign new_n701_ = \b[0]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] ) & (~\b[0]  | (~\a[11]  ^ ~\a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[1]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  ^ \a[14] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[0]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[1]  | (~\a[11]  ^ ~\a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[2]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  ^ \a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )));
  assign new_n702_ = \a[14]  ^ (((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[2]  | (~\a[11]  ^ ~\a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[3]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  ^ \a[14] )));
  assign new_n703_ = (\b[0]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) ^ ((~\b[0]  | (~\a[11]  ^ ~\a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[1]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  ^ \a[14] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[0]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[1]  | (~\a[11]  ^ ~\a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[2]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  ^ \a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n704_ = ((~\b[0]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  ^ ~\a[15] ) | (\a[15]  ^ \a[16] )) & (~\b[1]  | (~\a[14]  ^ ~\a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[2]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  ^ \a[17] )) & ((~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))) ^ (~\a[17]  | ((~\b[0]  | (~\a[14]  ^ ~\a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\b[1]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  ^ \a[17] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] )) & \a[17]  & (~\b[0]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ))));
  assign new_n705_ = ~new_n690_ ^ ((new_n613_ ^ ~new_n614_) ^ ((~new_n615_ & new_n623_) | (~new_n616_ & (new_n615_ | ~new_n623_) & (~new_n615_ | new_n623_))));
  assign new_n706_ = \a[14]  ^ (new_n707_ & (~new_n698_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n707_ = (~\b[8]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[9]  | (~\a[11]  ^ ~\a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[10]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  ^ \a[14] ));
  assign new_n708_ = \a[14]  ^ ((~\b[6]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[7]  | (\a[11]  ^ \a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[8]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  ^ \a[14] )) & ((\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n79_ & (~\b[7]  ^ \b[8] ))));
  assign new_n709_ = ~new_n685_ ^ (new_n610_ ^ ~new_n684_);
  assign new_n710_ = ~new_n682_ ^ (new_n624_ ^ ((~new_n627_ & (new_n471_ | (~new_n470_ & new_n478_) | (new_n470_ & ~new_n478_)) & (~new_n471_ | (~new_n470_ ^ new_n478_))) | (~new_n610_ & (new_n627_ | (~new_n471_ & (new_n470_ | ~new_n478_) & (~new_n470_ | new_n478_)) | (new_n471_ & (new_n470_ ^ new_n478_))) & (~new_n627_ | (~new_n471_ ^ (~new_n470_ ^ new_n478_))))));
  assign new_n711_ = \a[14]  ^ ((~\b[11]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[12]  | (\a[11]  ^ \a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[13]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  ^ \a[14] )) & (~new_n133_ | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n712_ = new_n677_ & (~new_n629_ ^ (new_n602_ | (~new_n605_ & new_n628_)));
  assign new_n713_ = \a[14]  ^ ((~\b[14]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[15]  | (\a[11]  ^ \a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[16]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  ^ \a[14] )) & (~new_n186_ | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n714_ = \a[14]  ^ ((~\b[12]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[13]  | (\a[11]  ^ \a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[14]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  ^ \a[14] )) & ((\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n142_ & (~\b[13]  ^ \b[14] ))));
  assign new_n715_ = ~new_n673_ ^ (new_n597_ ^ ~new_n672_);
  assign new_n716_ = ~new_n670_ ^ ((~new_n595_ & ~new_n631_) ^ ((~new_n633_ & (new_n460_ | ~new_n483_) & (~new_n460_ | new_n483_)) | (~new_n597_ & (new_n633_ | (~new_n460_ & new_n483_) | (new_n460_ & ~new_n483_)) & (~new_n633_ | (~new_n460_ ^ new_n483_)))));
  assign new_n717_ = \a[14]  ^ ((~\b[17]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[18]  | (\a[11]  ^ \a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[19]  | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  ^ \a[14] )) & (~new_n253_ | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n718_ = new_n665_ & (~new_n635_ ^ (new_n590_ | (~new_n593_ & new_n634_)));
  assign new_n719_ = \a[14]  ^ (((\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~new_n201_ ^ ~\b[19] )) & (~\b[18]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  ^ \a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[19]  | (\a[11]  ^ \a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )));
  assign new_n720_ = \a[14]  ^ (new_n577_ ^ ~new_n654_);
  assign new_n721_ = ((\a[11]  & (new_n643_ | (new_n642_ & \a[14] ) | (~new_n642_ & ~\a[14] )) & (~new_n643_ | (new_n642_ ^ \a[14] ))) | (((new_n723_ & \a[11] ) | (((new_n724_ & \a[11] ) | (~new_n725_ & (new_n724_ | \a[11] ) & (~new_n724_ | ~\a[11] ))) & (~new_n723_ | ~\a[11] ) & (new_n723_ | \a[11] ))) & (~\a[11]  | (~new_n643_ & (~new_n642_ | ~\a[14] ) & (new_n642_ | \a[14] )) | (new_n643_ & (~new_n642_ ^ \a[14] ))) & (\a[11]  | (~new_n643_ ^ (new_n642_ ^ \a[14] ))))) ^ (\a[11]  ^ (new_n722_ ^ ((new_n642_ & \a[14] ) | (~new_n643_ & (~new_n642_ | ~\a[14] ) & (new_n642_ | \a[14] )))));
  assign new_n722_ = \a[14]  ^ ((new_n562_ ^ \a[17] ) ^ ((new_n563_ & \a[17] ) | (~new_n564_ & (new_n563_ | \a[17] ) & (~new_n563_ | ~\a[17] ))));
  assign new_n723_ = ((\a[14]  & (new_n644_ | (new_n566_ & \a[17] ) | (~new_n566_ & ~\a[17] )) & (~new_n644_ | (new_n566_ ^ \a[17] ))) | (((new_n646_ & \a[14] ) | ((~new_n646_ | ~\a[14] ) & (new_n646_ | \a[14] ) & ((new_n647_ & \a[14] ) | (~new_n648_ & (~new_n647_ | ~\a[14] ) & (new_n647_ | \a[14] ))))) & (~\a[14]  | (~new_n644_ & (~new_n566_ | ~\a[17] ) & (new_n566_ | \a[17] )) | (new_n644_ & (~new_n566_ ^ \a[17] ))) & (\a[14]  | (~new_n644_ ^ (new_n566_ ^ \a[17] ))))) ^ (\a[14]  ^ (new_n645_ ^ ((new_n566_ & \a[17] ) | (~new_n644_ & (~new_n566_ | ~\a[17] ) & (new_n566_ | \a[17] )))));
  assign new_n724_ = ((new_n646_ & \a[14] ) | ((~new_n646_ | ~\a[14] ) & (new_n646_ | \a[14] ) & ((new_n647_ & \a[14] ) | (~new_n648_ & (new_n647_ | \a[14] ) & (~new_n647_ | ~\a[14] ))))) ^ (\a[14]  ^ (~new_n644_ ^ (~new_n566_ ^ ~\a[17] )));
  assign new_n725_ = (~\a[11]  | ((~new_n646_ | ~\a[14] ) & (new_n646_ | \a[14] ) & ((new_n647_ & \a[14] ) | ((~new_n647_ | ~\a[14] ) & (new_n647_ | \a[14] ) & ((new_n649_ & \a[14] ) | (~new_n726_ & (~new_n649_ | ~\a[14] ) & (new_n649_ | \a[14] )))))) | ((~new_n646_ ^ \a[14] ) & (~new_n647_ | ~\a[14] ) & ((new_n647_ & \a[14] ) | (~new_n647_ & ~\a[14] ) | ((~new_n649_ | ~\a[14] ) & (new_n726_ | (new_n649_ & \a[14] ) | (~new_n649_ & ~\a[14] )))))) & (((~\a[11]  | ((~new_n647_ | ~\a[14] ) & (new_n647_ | \a[14] ) & ((new_n649_ & \a[14] ) | (~new_n726_ & (~new_n649_ | ~\a[14] ) & (new_n649_ | \a[14] )))) | ((~new_n647_ ^ \a[14] ) & (~new_n649_ | ~\a[14] ) & (new_n726_ | (new_n649_ & \a[14] ) | (~new_n649_ & ~\a[14] )))) & (((~\a[11]  | (~new_n726_ & (~new_n649_ | ~\a[14] ) & (new_n649_ | \a[14] )) | (new_n726_ & (~new_n649_ ^ \a[14] ))) & (((~new_n727_ | ~\a[11] ) & (new_n728_ | (new_n727_ & \a[11] ) | (~new_n727_ & ~\a[11] ))) | (\a[11]  & (new_n726_ | (new_n649_ & \a[14] ) | (~new_n649_ & ~\a[14] )) & (~new_n726_ | (new_n649_ ^ \a[14] ))) | (~\a[11]  & (new_n726_ ^ (new_n649_ ^ \a[14] ))))) | (\a[11]  & ((new_n647_ & \a[14] ) | (~new_n647_ & ~\a[14] ) | ((~new_n649_ | ~\a[14] ) & (new_n726_ | (new_n649_ & \a[14] ) | (~new_n649_ & ~\a[14] )))) & ((new_n647_ ^ \a[14] ) | (new_n649_ & \a[14] ) | (~new_n726_ & (~new_n649_ | ~\a[14] ) & (new_n649_ | \a[14] )))) | (~\a[11]  & ((~new_n647_ ^ \a[14] ) ^ ((new_n649_ & \a[14] ) | (~new_n726_ & (~new_n649_ | ~\a[14] ) & (new_n649_ | \a[14] ))))))) | (\a[11]  & ((new_n646_ & \a[14] ) | (~new_n646_ & ~\a[14] ) | ((~new_n647_ | ~\a[14] ) & ((new_n647_ & \a[14] ) | (~new_n647_ & ~\a[14] ) | ((~new_n649_ | ~\a[14] ) & (new_n726_ | (new_n649_ & \a[14] ) | (~new_n649_ & ~\a[14] )))))) & ((new_n646_ ^ \a[14] ) | (new_n647_ & \a[14] ) | ((~new_n647_ | ~\a[14] ) & (new_n647_ | \a[14] ) & ((new_n649_ & \a[14] ) | (~new_n726_ & (~new_n649_ | ~\a[14] ) & (new_n649_ | \a[14] )))))) | (~\a[11]  & ((~new_n646_ ^ \a[14] ) ^ ((new_n647_ & \a[14] ) | ((~new_n647_ | ~\a[14] ) & (new_n647_ | \a[14] ) & ((new_n649_ & \a[14] ) | (~new_n726_ & (~new_n649_ | ~\a[14] ) & (new_n649_ | \a[14] ))))))));
  assign new_n726_ = (~\a[14]  | ((~new_n571_ | ~\a[17] ) & (new_n571_ | \a[17] ) & ((new_n572_ & \a[17] ) | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))))) | ((~new_n571_ ^ \a[17] ) & (~new_n572_ | ~\a[17] ) & ((new_n572_ & \a[17] ) | (~new_n572_ & ~\a[17] ) | ((~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))))) & ((\a[14]  & ((new_n571_ & \a[17] ) | (~new_n571_ & ~\a[17] ) | ((~new_n572_ | ~\a[17] ) & ((new_n572_ & \a[17] ) | (~new_n572_ & ~\a[17] ) | ((~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))))) & ((new_n571_ ^ \a[17] ) | (new_n572_ & \a[17] ) | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))))) | (~\a[14]  & ((~new_n571_ ^ \a[17] ) ^ ((new_n572_ & \a[17] ) | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] ))))))) | ((~\a[14]  | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))) | ((~new_n572_ ^ \a[17] ) & (~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))) & ((\a[14]  & ((new_n572_ & \a[17] ) | (~new_n572_ & ~\a[17] ) | ((~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))) & ((new_n572_ ^ \a[17] ) | (new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))) | (~\a[14]  & ((~new_n572_ ^ \a[17] ) ^ ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] ))))) | ((~\a[14]  | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )) | (new_n575_ & (~new_n573_ ^ \a[17] ))) & (new_n650_ | (\a[14]  & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )) & (~new_n575_ | (new_n573_ ^ \a[17] ))) | (~\a[14]  & (new_n575_ ^ (new_n573_ ^ \a[17] ))))))));
  assign new_n727_ = (\a[14]  ^ ((new_n571_ ^ \a[17] ) ^ ((new_n572_ & \a[17] ) | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] ))))))) ^ ((\a[14]  & ((new_n572_ & \a[17] ) | (~new_n572_ & ~\a[17] ) | ((~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))) & ((new_n572_ ^ \a[17] ) | (new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))) | ((~\a[14]  | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))) | ((~new_n572_ ^ \a[17] ) & (~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))) & (\a[14]  | ((new_n572_ ^ \a[17] ) ^ ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] ))))) & ((\a[14]  & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )) & (~new_n575_ | (new_n573_ ^ \a[17] ))) | (~new_n650_ & (~\a[14]  | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )) | (new_n575_ & (~new_n573_ ^ \a[17] ))) & (\a[14]  | (~new_n575_ ^ (new_n573_ ^ \a[17] )))))));
  assign new_n728_ = (~\a[11]  | (new_n729_ & ~new_n731_) | (~new_n729_ & new_n731_)) & ((\a[11]  & (~new_n729_ | new_n731_) & (new_n729_ | ~new_n731_)) | (~\a[11]  & (~new_n729_ ^ ~new_n731_)) | ((~new_n732_ | ~\a[11] ) & ((new_n732_ & \a[11] ) | (~new_n732_ & ~\a[11] ) | ((~new_n733_ | ~\a[11] ) & ((new_n733_ & \a[11] ) | (~new_n733_ & ~\a[11] ) | (~new_n734_ & (new_n735_ | ~new_n806_)))))));
  assign new_n729_ = (~\a[14]  | (new_n575_ & ~new_n730_) | (~new_n575_ & new_n730_)) & ((\a[14]  & (~new_n575_ | new_n730_) & (new_n575_ | ~new_n730_)) | (~\a[14]  & (~new_n575_ ^ ~new_n730_)) | ((~new_n651_ | ~\a[14] ) & ((new_n651_ & \a[14] ) | (~new_n651_ & ~\a[14] ) | ((~new_n652_ | ~\a[14] ) & ((new_n652_ & \a[14] ) | (~new_n652_ & ~\a[14] ) | (~new_n653_ & (new_n655_ | ~new_n720_)))))));
  assign new_n730_ = \a[17]  ^ (new_n431_ ^ ~new_n574_);
  assign new_n731_ = \a[14]  ^ ((new_n572_ ^ \a[17] ) ^ ((new_n573_ & \a[17] ) | (~new_n575_ & (new_n573_ | \a[17] ) & (~new_n573_ | ~\a[17] ))));
  assign new_n732_ = (\a[14]  ^ (new_n575_ ^ ~new_n730_)) ^ ((new_n651_ & \a[14] ) | ((~new_n651_ | ~\a[14] ) & (new_n651_ | \a[14] ) & ((new_n652_ & \a[14] ) | ((~new_n652_ | ~\a[14] ) & (new_n652_ | \a[14] ) & (new_n653_ | (~new_n655_ & new_n720_))))));
  assign new_n733_ = (new_n651_ ^ \a[14] ) ^ ((new_n652_ & \a[14] ) | ((~new_n652_ | ~\a[14] ) & (new_n652_ | \a[14] ) & (new_n653_ | (~new_n655_ & new_n720_))));
  assign new_n734_ = \a[11]  & ((new_n652_ & \a[14] ) | (~new_n652_ & ~\a[14] ) | (~new_n653_ & (new_n655_ | ~new_n720_))) & ((new_n652_ ^ \a[14] ) | new_n653_ | (~new_n655_ & new_n720_));
  assign new_n735_ = (~\a[11]  | (new_n655_ & ~new_n720_) | (~new_n655_ & new_n720_)) & ((\a[11]  & (~new_n655_ | new_n720_) & (new_n655_ | ~new_n720_)) | (~\a[11]  & (~new_n655_ ^ ~new_n720_)) | ((~new_n736_ | ~\a[11] ) & ((new_n736_ & \a[11] ) | (~new_n736_ & ~\a[11] ) | ((~new_n737_ | ~\a[11] ) & ((new_n737_ & \a[11] ) | (~new_n737_ & ~\a[11] ) | (~new_n738_ & (new_n740_ | ~new_n805_)))))));
  assign new_n736_ = (new_n657_ ^ \a[14] ) ^ ((\a[14]  & ((new_n656_ & \a[17] ) | (~new_n656_ & ~\a[17] ) | ((~new_n579_ | ~\a[17] ) & ((new_n579_ & \a[17] ) | (~new_n579_ & ~\a[17] ) | ((~new_n580_ | ~\a[17] ) & (new_n581_ | (new_n580_ & \a[17] ) | (~new_n580_ & ~\a[17] )))))) & ((new_n656_ ^ \a[17] ) | (new_n579_ & \a[17] ) | ((~new_n579_ | ~\a[17] ) & (new_n579_ | \a[17] ) & ((new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] )))))) | ((~\a[14]  | ((~new_n656_ | ~\a[17] ) & (new_n656_ | \a[17] ) & ((new_n579_ & \a[17] ) | ((~new_n579_ | ~\a[17] ) & (new_n579_ | \a[17] ) & ((new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] )))))) | ((~new_n656_ ^ \a[17] ) & (~new_n579_ | ~\a[17] ) & ((new_n579_ & \a[17] ) | (~new_n579_ & ~\a[17] ) | ((~new_n580_ | ~\a[17] ) & (new_n581_ | (new_n580_ & \a[17] ) | (~new_n580_ & ~\a[17] )))))) & (\a[14]  | ((new_n656_ ^ \a[17] ) ^ ((new_n579_ & \a[17] ) | ((~new_n579_ | ~\a[17] ) & (new_n579_ | \a[17] ) & ((new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] ))))))) & ((\a[14]  & ((new_n579_ & \a[17] ) | (~new_n579_ & ~\a[17] ) | ((~new_n580_ | ~\a[17] ) & (new_n581_ | (new_n580_ & \a[17] ) | (~new_n580_ & ~\a[17] )))) & ((new_n579_ ^ \a[17] ) | (new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] )))) | (~new_n658_ & (~\a[14]  | ((~new_n579_ | ~\a[17] ) & (new_n579_ | \a[17] ) & ((new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] )))) | ((~new_n579_ ^ \a[17] ) & (~new_n580_ | ~\a[17] ) & (new_n581_ | (new_n580_ & \a[17] ) | (~new_n580_ & ~\a[17] )))) & (\a[14]  | ((new_n579_ ^ \a[17] ) ^ ((new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] )))))))));
  assign new_n737_ = (\a[14]  ^ ((~new_n656_ ^ ~\a[17] ) ^ ((new_n579_ & \a[17] ) | ((~new_n579_ | ~\a[17] ) & (new_n579_ | \a[17] ) & ((new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] ))))))) ^ ((\a[14]  & ((new_n579_ & \a[17] ) | (~new_n579_ & ~\a[17] ) | ((~new_n580_ | ~\a[17] ) & (new_n581_ | (new_n580_ & \a[17] ) | (~new_n580_ & ~\a[17] )))) & ((new_n579_ ^ \a[17] ) | (new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] )))) | (~new_n658_ & (~\a[14]  | ((~new_n579_ | ~\a[17] ) & (new_n579_ | \a[17] ) & ((new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] )))) | ((~new_n579_ ^ \a[17] ) & (~new_n580_ | ~\a[17] ) & (new_n581_ | (new_n580_ & \a[17] ) | (~new_n580_ & ~\a[17] )))) & (\a[14]  | ((new_n579_ ^ \a[17] ) ^ ((new_n580_ & \a[17] ) | (~new_n581_ & (~new_n580_ | ~\a[17] ) & (new_n580_ | \a[17] )))))));
  assign new_n738_ = \a[11]  & (~new_n658_ | new_n739_) & (new_n658_ | ~new_n739_);
  assign new_n739_ = \a[14]  ^ ((new_n579_ ^ \a[17] ) ^ ((new_n580_ & \a[17] ) | (~new_n581_ & (new_n580_ | \a[17] ) & (~new_n580_ | ~\a[17] ))));
  assign new_n740_ = (~new_n742_ | ~\a[11] ) & ((new_n742_ & \a[11] ) | (~new_n742_ & ~\a[11] ) | ((~\a[11]  | ((~new_n741_ | ~\a[14] ) & (new_n741_ | \a[14] ) & ((~new_n660_ & \a[14] ) | (((new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] ))) & (new_n660_ | ~\a[14] ) & (~new_n660_ | \a[14] )))) | ((~new_n741_ ^ \a[14] ) & (new_n660_ | ~\a[14] ) & (((~new_n661_ | ~\a[14] ) & (new_n662_ | (new_n661_ & \a[14] ) | (~new_n661_ & ~\a[14] ))) | (~new_n660_ & \a[14] ) | (new_n660_ & ~\a[14] )))) & (((~\a[11]  | (((new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] ))) & (new_n660_ | ~\a[14] ) & (~new_n660_ | \a[14] )) | ((~new_n661_ | ~\a[14] ) & (new_n662_ | (new_n661_ & \a[14] ) | (~new_n661_ & ~\a[14] )) & (new_n660_ ^ \a[14] ))) & (new_n743_ | (\a[11]  & (((~new_n661_ | ~\a[14] ) & (new_n662_ | (new_n661_ & \a[14] ) | (~new_n661_ & ~\a[14] ))) | (~new_n660_ & \a[14] ) | (new_n660_ & ~\a[14] )) & ((new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] )) | (~new_n660_ ^ \a[14] ))) | (~\a[11]  & (((~new_n661_ | ~\a[14] ) & (new_n662_ | (new_n661_ & \a[14] ) | (~new_n661_ & ~\a[14] ))) ^ (~new_n660_ ^ \a[14] ))))) | (\a[11]  & ((new_n741_ & \a[14] ) | (~new_n741_ & ~\a[14] ) | ((new_n660_ | ~\a[14] ) & (((~new_n661_ | ~\a[14] ) & (new_n662_ | (new_n661_ & \a[14] ) | (~new_n661_ & ~\a[14] ))) | (~new_n660_ & \a[14] ) | (new_n660_ & ~\a[14] )))) & ((new_n741_ ^ \a[14] ) | (~new_n660_ & \a[14] ) | (((new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] ))) & (new_n660_ | ~\a[14] ) & (~new_n660_ | \a[14] )))) | (~\a[11]  & ((~new_n741_ ^ \a[14] ) ^ ((~new_n660_ & \a[14] ) | (((new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] ))) & (new_n660_ | ~\a[14] ) & (~new_n660_ | \a[14] ))))))));
  assign new_n741_ = ~new_n659_ ^ (new_n582_ ^ \a[17] );
  assign new_n742_ = (\a[14]  ^ ((new_n580_ ^ \a[17] ) ^ ((new_n582_ & \a[17] ) | (~new_n659_ & (~new_n582_ | ~\a[17] ) & (new_n582_ | \a[17] ))))) ^ ((\a[14]  & (new_n659_ | (new_n582_ & \a[17] ) | (~new_n582_ & ~\a[17] )) & (~new_n659_ | (new_n582_ ^ \a[17] ))) | ((~\a[14]  | (~new_n659_ & (~new_n582_ | ~\a[17] ) & (new_n582_ | \a[17] )) | (new_n659_ & (~new_n582_ ^ \a[17] ))) & (\a[14]  | (~new_n659_ ^ (new_n582_ ^ \a[17] ))) & ((~new_n660_ & \a[14] ) | ((new_n660_ | ~\a[14] ) & (~new_n660_ | \a[14] ) & ((new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] )))))));
  assign new_n743_ = (~\a[11]  | ((~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] ) & ((new_n663_ & \a[14] ) | (~new_n744_ & (~new_n663_ | ~\a[14] ) & (new_n663_ | \a[14] )))) | ((~new_n661_ ^ \a[14] ) & (~new_n663_ | ~\a[14] ) & (new_n744_ | (new_n663_ & \a[14] ) | (~new_n663_ & ~\a[14] )))) & ((\a[11]  & ((new_n661_ & \a[14] ) | (~new_n661_ & ~\a[14] ) | ((~new_n663_ | ~\a[14] ) & (new_n744_ | (new_n663_ & \a[14] ) | (~new_n663_ & ~\a[14] )))) & ((new_n661_ ^ \a[14] ) | (new_n663_ & \a[14] ) | (~new_n744_ & (~new_n663_ | ~\a[14] ) & (new_n663_ | \a[14] )))) | (~\a[11]  & ((~new_n661_ ^ \a[14] ) ^ ((new_n663_ & \a[14] ) | (~new_n744_ & (~new_n663_ | ~\a[14] ) & (new_n663_ | \a[14] ))))) | ((~\a[11]  | (~new_n744_ & (~new_n663_ | ~\a[14] ) & (new_n663_ | \a[14] )) | (new_n744_ & (~new_n663_ ^ \a[14] ))) & ((\a[11]  & (new_n744_ | (new_n663_ & \a[14] ) | (~new_n663_ & ~\a[14] )) & (~new_n744_ | (new_n663_ ^ \a[14] ))) | (~\a[11]  & (new_n744_ ^ (new_n663_ ^ \a[14] ))) | ((new_n745_ | ~\a[11] ) & ((~new_n745_ & \a[11] ) | (new_n745_ & ~\a[11] ) | ((~new_n746_ | ~\a[11] ) & (new_n747_ | (new_n746_ & \a[11] ) | (~new_n746_ & ~\a[11] ))))))));
  assign new_n744_ = ~new_n664_ & (new_n718_ | ((new_n719_ | (~new_n593_ & new_n634_) | (new_n593_ & ~new_n634_)) & (new_n666_ | (~new_n719_ & (new_n593_ | ~new_n634_) & (~new_n593_ | new_n634_)) | (new_n719_ & (new_n593_ ^ new_n634_)))));
  assign new_n745_ = (~new_n664_ & ~new_n718_) ^ ((new_n719_ | (~new_n593_ & new_n634_) | (new_n593_ & ~new_n634_)) & (new_n666_ | (~new_n719_ & (new_n593_ | ~new_n634_) & (~new_n593_ | new_n634_)) | (new_n719_ & (new_n593_ ^ new_n634_))));
  assign new_n746_ = ~new_n666_ ^ (~new_n719_ ^ (~new_n593_ ^ new_n634_));
  assign new_n747_ = (~new_n748_ | ~\a[11] ) & ((new_n748_ & \a[11] ) | (~new_n748_ & ~\a[11] ) | (~new_n749_ & (new_n749_ | new_n803_ | ((new_n804_ | (~new_n674_ & new_n715_) | (new_n674_ & ~new_n715_)) & (new_n751_ | (~new_n804_ & (new_n674_ | ~new_n715_) & (~new_n674_ | new_n715_)) | (new_n804_ & (new_n674_ ^ new_n715_)))))));
  assign new_n748_ = (new_n667_ ^ ~new_n717_) ^ (new_n669_ | (new_n716_ & (new_n671_ | (~new_n674_ & new_n715_))));
  assign new_n749_ = ~new_n750_ & (~new_n716_ | (~new_n671_ & (new_n674_ | ~new_n715_))) & (new_n716_ | new_n671_ | (~new_n674_ & new_n715_));
  assign new_n750_ = \a[11]  ^ (~\b[19]  | (((\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (new_n201_ | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ))));
  assign new_n751_ = (~new_n752_ | new_n802_) & ((new_n752_ & ~new_n802_) | (~new_n752_ & new_n802_) | (~new_n754_ & (~new_n801_ | (~new_n756_ & (new_n759_ | ~new_n800_)))));
  assign new_n752_ = new_n753_ ^ (new_n676_ | (((~new_n714_ & (new_n605_ | ~new_n628_) & (~new_n605_ | new_n628_)) | (~new_n678_ & (new_n714_ | (~new_n605_ & new_n628_) | (new_n605_ & ~new_n628_)) & (~new_n714_ | (~new_n605_ ^ new_n628_)))) & ~new_n676_ & ~new_n712_));
  assign new_n753_ = ~new_n713_ ^ ((new_n600_ | (new_n629_ & (new_n602_ | (~new_n605_ & new_n628_)))) ^ (new_n598_ ^ ~new_n630_));
  assign new_n754_ = ~new_n755_ & (new_n676_ | new_n712_ | ((new_n714_ | (~new_n605_ & new_n628_) | (new_n605_ & ~new_n628_)) & (new_n678_ | (~new_n714_ & (new_n605_ | ~new_n628_) & (~new_n605_ | new_n628_)) | (new_n714_ & (new_n605_ ^ new_n628_))))) & ((~new_n676_ & ~new_n712_) | (~new_n714_ & (new_n605_ | ~new_n628_) & (~new_n605_ | new_n628_)) | (~new_n678_ & (new_n714_ | (~new_n605_ & new_n628_) | (new_n605_ & ~new_n628_)) & (~new_n714_ | (~new_n605_ ^ new_n628_))));
  assign new_n755_ = \a[11]  ^ ((~new_n199_ | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[17]  | (\a[8]  ^ \a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[18]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[16]  | (\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n756_ = ~new_n758_ & (~new_n678_ | new_n757_) & (new_n678_ | ~new_n757_);
  assign new_n757_ = ~new_n714_ ^ (new_n605_ ^ ~new_n628_);
  assign new_n758_ = \a[11]  ^ ((~new_n144_ | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[16]  | (\a[8]  ^ \a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[17]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[15]  | (\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n759_ = (~new_n760_ | new_n798_) & ((new_n760_ & ~new_n798_) | (~new_n760_ & new_n798_) | (~new_n761_ & (new_n761_ | new_n797_ | ((new_n799_ | (~new_n686_ & new_n709_) | (new_n686_ & ~new_n709_)) & (new_n763_ | (~new_n799_ & (new_n686_ | ~new_n709_) & (~new_n686_ | new_n709_)) | (new_n799_ & (new_n686_ ^ new_n709_)))))));
  assign new_n760_ = (new_n679_ ^ ~new_n711_) ^ (new_n681_ | (new_n710_ & (new_n683_ | (~new_n686_ & new_n709_))));
  assign new_n761_ = ~new_n762_ & (~new_n710_ | (~new_n683_ & (new_n686_ | ~new_n709_))) & (new_n710_ | new_n683_ | (~new_n686_ & new_n709_));
  assign new_n762_ = \a[11]  ^ ((((~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] ) & ((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )))) | ((~\b[14]  ^ \b[15] ) & (~\b[13]  | ~\b[14] ) & (new_n142_ | (\b[13]  & \b[14] ) | (~\b[13]  & ~\b[14] ))) | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[14]  | (\a[8]  ^ \a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[15]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[13]  | (\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n763_ = (~new_n764_ | new_n796_) & ((new_n764_ & ~new_n796_) | (~new_n764_ & new_n796_) | (~new_n766_ & (~new_n795_ | (~new_n768_ & (new_n771_ | ~new_n794_)))));
  assign new_n764_ = new_n765_ ^ (new_n689_ | (new_n705_ & ((~new_n708_ & (new_n616_ | (~new_n615_ & new_n623_) | (new_n615_ & ~new_n623_)) & (~new_n616_ | (~new_n615_ ^ new_n623_))) | (~new_n691_ & (new_n708_ | (~new_n616_ & (new_n615_ | ~new_n623_) & (~new_n615_ | new_n623_)) | (new_n616_ & (new_n615_ ^ new_n623_))) & (~new_n708_ | (~new_n616_ ^ (~new_n615_ ^ new_n623_)))))));
  assign new_n765_ = ~new_n706_ ^ ((new_n611_ ^ ~new_n612_) ^ ((new_n613_ & ~new_n614_) | ((~new_n613_ | new_n614_) & (new_n613_ | ~new_n614_) & ((~new_n615_ & new_n623_) | (~new_n616_ & (new_n615_ | ~new_n623_) & (~new_n615_ | new_n623_))))));
  assign new_n766_ = ~new_n767_ & (~new_n705_ | ((new_n708_ | (~new_n616_ & (new_n615_ | ~new_n623_) & (~new_n615_ | new_n623_)) | (new_n616_ & (new_n615_ ^ new_n623_))) & (new_n691_ | (~new_n708_ & (new_n616_ | (~new_n615_ & new_n623_) | (new_n615_ & ~new_n623_)) & (~new_n616_ | (~new_n615_ ^ new_n623_))) | (new_n708_ & (new_n616_ ^ (~new_n615_ ^ new_n623_)))))) & (new_n705_ | (~new_n708_ & (new_n616_ | (~new_n615_ & new_n623_) | (new_n615_ & ~new_n623_)) & (~new_n616_ | (~new_n615_ ^ new_n623_))) | (~new_n691_ & (new_n708_ | (~new_n616_ & (new_n615_ | ~new_n623_) & (~new_n615_ | new_n623_)) | (new_n616_ & (new_n615_ ^ new_n623_))) & (~new_n708_ | (~new_n616_ ^ (~new_n615_ ^ new_n623_)))));
  assign new_n767_ = \a[11]  ^ ((~new_n107_ | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[11]  | (\a[8]  ^ \a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[12]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[10]  | (\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n768_ = ~new_n770_ & (~new_n691_ | new_n769_) & (new_n691_ | ~new_n769_);
  assign new_n769_ = ~new_n708_ ^ (~new_n616_ ^ (~new_n615_ ^ new_n623_));
  assign new_n770_ = \a[11]  ^ ((~new_n135_ | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[10]  | (\a[8]  ^ \a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[11]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[9]  | (\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n771_ = (~new_n773_ | new_n791_) & ((~new_n774_ & (~new_n790_ | ((new_n793_ | (new_n772_ & ~new_n697_) | (~new_n772_ & new_n697_)) & (new_n776_ | (~new_n793_ & (~new_n772_ | new_n697_) & (new_n772_ | ~new_n697_)) | (new_n793_ & (~new_n772_ ^ ~new_n697_)))))) | (new_n773_ & ~new_n791_) | (~new_n773_ & new_n791_));
  assign new_n772_ = new_n696_ ^ ~new_n704_;
  assign new_n773_ = (new_n692_ ^ ~new_n693_) ^ ((new_n694_ & ~new_n695_) | (((~new_n696_ & new_n704_) | (~new_n697_ & (new_n696_ | ~new_n704_) & (~new_n696_ | new_n704_))) & (~new_n694_ | new_n695_) & (new_n694_ | ~new_n695_)));
  assign new_n774_ = ~new_n775_ & ((new_n694_ & ~new_n695_) | (~new_n694_ & new_n695_) | ((new_n696_ | ~new_n704_) & (new_n697_ | (~new_n696_ & new_n704_) | (new_n696_ & ~new_n704_)))) & ((new_n694_ ^ ~new_n695_) | (~new_n696_ & new_n704_) | (~new_n697_ & (new_n696_ | ~new_n704_) & (~new_n696_ | new_n704_)));
  assign new_n775_ = \a[11]  ^ ((((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))) | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[8]  | (\a[8]  ^ \a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[9]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[7]  | (\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n776_ = (new_n777_ | ~new_n778_) & ((new_n777_ & ~new_n778_) | (~new_n777_ & new_n778_) | ((~new_n779_ | new_n780_) & (((new_n781_ | ~new_n789_) & (new_n782_ | (~new_n781_ & new_n789_) | (new_n781_ & ~new_n789_))) | (new_n779_ & ~new_n780_) | (~new_n779_ & new_n780_))));
  assign new_n777_ = \a[11]  ^ ((~new_n88_ | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[6]  | (\a[8]  ^ \a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[7]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[5]  | (\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n778_ = (new_n701_ | (~new_n702_ & new_n703_)) ^ (new_n700_ ^ (~\a[14]  ^ (new_n699_ & (~new_n98_ | ~new_n698_))));
  assign new_n779_ = new_n702_ ^ ~new_n703_;
  assign new_n780_ = \a[11]  ^ ((~new_n91_ | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[5]  | (\a[8]  ^ \a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[6]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[4]  | (\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n781_ = \a[11]  ^ ((~new_n94_ | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[4]  | (\a[8]  ^ \a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[5]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[3]  | (\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n782_ = (~new_n785_ | (\a[11]  ^ (new_n784_ & (~new_n98_ | ~new_n783_)))) & ((~new_n786_ & (new_n787_ | ~new_n788_)) | (new_n785_ & (~\a[11]  ^ (new_n784_ & (~new_n98_ | ~new_n783_)))) | (~new_n785_ & (~\a[11]  | ~new_n784_ | (new_n98_ & new_n783_)) & (\a[11]  | (new_n784_ & (~new_n98_ | ~new_n783_)))));
  assign new_n783_ = (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (~\a[10]  | ~\a[11] ) & (\a[10]  | \a[11] );
  assign new_n784_ = (~\b[3]  | (~\a[8]  ^ ~\a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[4]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[2]  | (\a[9]  ^ \a[10] ) | (~\a[8]  ^ ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ));
  assign new_n785_ = ((\b[0]  & (\a[11]  ^ ~\a[12] ) & (~\a[12]  | ~\a[13] ) & (\a[12]  | \a[13] )) | (\b[1]  & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ) & (~\a[13]  ^ \a[14] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ) & (~\a[13]  | ~\a[14] ) & (\a[13]  | \a[14] ))) ^ (\a[14]  & \b[0]  & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ));
  assign new_n786_ = \b[0]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] ) & (~\b[0]  | (~\a[8]  ^ ~\a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[1]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  ^ \a[11] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[0]  | (\a[9]  ^ \a[10] ) | (~\a[8]  ^ ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[1]  | (~\a[8]  ^ ~\a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[2]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  ^ \a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )));
  assign new_n787_ = \a[11]  ^ (((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (~\a[8]  ^ ~\a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[3]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[1]  | (\a[9]  ^ \a[10] ) | (~\a[8]  ^ ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n788_ = (\b[0]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] )) ^ ((~\b[0]  | (~\a[8]  ^ ~\a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[1]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  ^ \a[11] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[0]  | (\a[9]  ^ \a[10] ) | (~\a[8]  ^ ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[1]  | (~\a[8]  ^ ~\a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[2]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  ^ \a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n789_ = ((~\b[0]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  ^ ~\a[12] ) | (\a[12]  ^ \a[13] )) & (~\b[1]  | (~\a[11]  ^ ~\a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[2]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  ^ \a[14] )) & ((~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))) ^ (~\a[14]  | ((~\b[0]  | (~\a[11]  ^ ~\a[12] ) | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] )) & (~\b[1]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  ^ \a[14] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ))));
  assign new_n790_ = ~new_n775_ ^ ((new_n694_ ^ ~new_n695_) ^ ((~new_n696_ & new_n704_) | (~new_n697_ & (new_n696_ | ~new_n704_) & (~new_n696_ | new_n704_))));
  assign new_n791_ = \a[11]  ^ (new_n792_ & (~new_n783_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n792_ = (~\b[9]  | (~\a[8]  ^ ~\a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[10]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[8]  | (\a[9]  ^ \a[10] ) | (~\a[8]  ^ ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ));
  assign new_n793_ = \a[11]  ^ ((~\b[7]  | (\a[8]  ^ \a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[8]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[6]  | (\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & ((\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n79_ & (~\b[7]  ^ \b[8] ))));
  assign new_n794_ = ~new_n770_ ^ (new_n691_ ^ ~new_n769_);
  assign new_n795_ = ~new_n767_ ^ (new_n705_ ^ ((~new_n708_ & (new_n616_ | (~new_n615_ & new_n623_) | (new_n615_ & ~new_n623_)) & (~new_n616_ | (~new_n615_ ^ new_n623_))) | (~new_n691_ & (new_n708_ | (~new_n616_ & (new_n615_ | ~new_n623_) & (~new_n615_ | new_n623_)) | (new_n616_ & (new_n615_ ^ new_n623_))) & (~new_n708_ | (~new_n616_ ^ (~new_n615_ ^ new_n623_))))));
  assign new_n796_ = \a[11]  ^ ((~new_n133_ | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[12]  | (\a[8]  ^ \a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[13]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[11]  | (\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n797_ = new_n762_ & (~new_n710_ ^ (new_n683_ | (~new_n686_ & new_n709_)));
  assign new_n798_ = \a[11]  ^ ((~new_n186_ | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[15]  | (\a[8]  ^ \a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[16]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[14]  | (\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n799_ = \a[11]  ^ ((~\b[13]  | (\a[8]  ^ \a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[14]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[12]  | (\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & ((\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n142_ & (~\b[13]  ^ \b[14] ))));
  assign new_n800_ = ~new_n758_ ^ (new_n678_ ^ ~new_n757_);
  assign new_n801_ = ~new_n755_ ^ ((~new_n676_ & ~new_n712_) ^ ((~new_n714_ & (new_n605_ | ~new_n628_) & (~new_n605_ | new_n628_)) | (~new_n678_ & (new_n714_ | (~new_n605_ & new_n628_) | (new_n605_ & ~new_n628_)) & (~new_n714_ | (~new_n605_ ^ new_n628_)))));
  assign new_n802_ = \a[11]  ^ ((~new_n253_ | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & (~\b[18]  | (\a[8]  ^ \a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[19]  | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  ^ \a[11] )) & (~\b[17]  | (\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n803_ = new_n750_ & (~new_n716_ ^ (new_n671_ | (~new_n674_ & new_n715_)));
  assign new_n804_ = \a[11]  ^ (((\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~new_n201_ ^ ~\b[19] )) & (~\b[19]  | (\a[8]  ^ \a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[18]  | (\a[9]  ^ \a[10] ) | (\a[8]  ^ \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n805_ = \a[11]  ^ (new_n658_ ^ ~new_n739_);
  assign new_n806_ = \a[11]  ^ ((new_n652_ ^ \a[14] ) ^ (new_n653_ | (~new_n655_ & new_n720_)));
  assign new_n807_ = (~new_n808_ | ~\a[8] ) & ((~new_n808_ & ~\a[8] ) | (new_n808_ & \a[8] ) | ((~new_n809_ | ~\a[8] ) & ((new_n809_ & \a[8] ) | (~new_n809_ & ~\a[8] ) | ((~\a[8]  | ((~new_n893_ | ~\a[11] ) & (new_n893_ | \a[11] ) & ((new_n727_ & \a[11] ) | (~new_n728_ & (~new_n727_ | ~\a[11] ) & (new_n727_ | \a[11] )))) | ((~new_n893_ ^ \a[11] ) & (~new_n727_ | ~\a[11] ) & (new_n728_ | (new_n727_ & \a[11] ) | (~new_n727_ & ~\a[11] )))) & (new_n810_ | (\a[8]  & ((new_n893_ & \a[11] ) | (~new_n893_ & ~\a[11] ) | ((~new_n727_ | ~\a[11] ) & (new_n728_ | (new_n727_ & \a[11] ) | (~new_n727_ & ~\a[11] )))) & ((new_n893_ ^ \a[11] ) | (new_n727_ & \a[11] ) | (~new_n728_ & (~new_n727_ | ~\a[11] ) & (new_n727_ | \a[11] )))) | (~\a[8]  & ((~new_n893_ ^ \a[11] ) ^ ((new_n727_ & \a[11] ) | (~new_n728_ & (~new_n727_ | ~\a[11] ) & (new_n727_ | \a[11] ))))))))));
  assign new_n808_ = ((\a[11]  & ((new_n647_ & \a[14] ) | (~new_n647_ & ~\a[14] ) | ((~new_n649_ | ~\a[14] ) & (new_n726_ | (new_n649_ & \a[14] ) | (~new_n649_ & ~\a[14] )))) & ((new_n647_ ^ \a[14] ) | (new_n649_ & \a[14] ) | (~new_n726_ & (~new_n649_ | ~\a[14] ) & (new_n649_ | \a[14] )))) | (((\a[11]  & (new_n726_ | (new_n649_ & \a[14] ) | (~new_n649_ & ~\a[14] )) & (~new_n726_ | (new_n649_ ^ \a[14] ))) | (((new_n727_ & \a[11] ) | (~new_n728_ & (~new_n727_ | ~\a[11] ) & (new_n727_ | \a[11] ))) & (~\a[11]  | (~new_n726_ & (~new_n649_ | ~\a[14] ) & (new_n649_ | \a[14] )) | (new_n726_ & (~new_n649_ ^ \a[14] ))) & (\a[11]  | (~new_n726_ ^ (new_n649_ ^ \a[14] ))))) & (~\a[11]  | ((~new_n647_ | ~\a[14] ) & (new_n647_ | \a[14] ) & ((new_n649_ & \a[14] ) | (~new_n726_ & (~new_n649_ | ~\a[14] ) & (new_n649_ | \a[14] )))) | ((~new_n647_ ^ \a[14] ) & (~new_n649_ | ~\a[14] ) & (new_n726_ | (new_n649_ & \a[14] ) | (~new_n649_ & ~\a[14] )))) & (\a[11]  | ((new_n647_ ^ \a[14] ) ^ ((new_n649_ & \a[14] ) | (~new_n726_ & (~new_n649_ | ~\a[14] ) & (new_n649_ | \a[14] ))))))) ^ (\a[11]  ^ ((new_n646_ ^ \a[14] ) ^ ((new_n647_ & \a[14] ) | ((~new_n647_ | ~\a[14] ) & (new_n647_ | \a[14] ) & ((new_n649_ & \a[14] ) | (~new_n726_ & (~new_n649_ | ~\a[14] ) & (new_n649_ | \a[14] )))))));
  assign new_n809_ = ((\a[11]  & (new_n726_ | (~new_n649_ & ~\a[14] ) | (new_n649_ & \a[14] )) & (~new_n726_ | (~new_n649_ ^ ~\a[14] ))) | (((new_n727_ & \a[11] ) | (~new_n728_ & (new_n727_ | \a[11] ) & (~new_n727_ | ~\a[11] ))) & (~\a[11]  | (~new_n726_ & (new_n649_ | \a[14] ) & (~new_n649_ | ~\a[14] )) | (new_n726_ & (new_n649_ ^ ~\a[14] ))) & (\a[11]  | (~new_n726_ ^ (~new_n649_ ^ ~\a[14] ))))) ^ (\a[11]  ^ ((~new_n647_ ^ ~\a[14] ) ^ ((new_n649_ & \a[14] ) | (~new_n726_ & (new_n649_ | \a[14] ) & (~new_n649_ | ~\a[14] )))));
  assign new_n810_ = (~\a[8]  | (new_n814_ & (new_n811_ | (~new_n812_ & new_n813_))) | (~new_n814_ & ~new_n811_ & (new_n812_ | ~new_n813_))) & (((~\a[8]  | (~new_n812_ & new_n813_) | (new_n812_ & ~new_n813_)) & (((~new_n815_ | ~\a[8] ) & ((new_n815_ & \a[8] ) | (~new_n815_ & ~\a[8] ) | ((~new_n816_ | ~\a[8] ) & (new_n817_ | (new_n816_ & \a[8] ) | (~new_n816_ & ~\a[8] ))))) | (\a[8]  & (new_n812_ | ~new_n813_) & (~new_n812_ | new_n813_)) | (~\a[8]  & (new_n812_ ^ new_n813_)))) | (\a[8]  & (~new_n814_ | (~new_n811_ & (new_n812_ | ~new_n813_))) & (new_n814_ | new_n811_ | (~new_n812_ & new_n813_))) | (~\a[8]  & (~new_n814_ ^ (new_n811_ | (~new_n812_ & new_n813_)))));
  assign new_n811_ = \a[11]  & (~new_n729_ | new_n731_) & (new_n729_ | ~new_n731_);
  assign new_n812_ = (~new_n732_ | ~\a[11] ) & ((new_n732_ & \a[11] ) | (~new_n732_ & ~\a[11] ) | ((~new_n733_ | ~\a[11] ) & ((new_n733_ & \a[11] ) | (~new_n733_ & ~\a[11] ) | (~new_n734_ & (new_n735_ | ~new_n806_)))));
  assign new_n813_ = \a[11]  ^ (new_n729_ ^ ~new_n731_);
  assign new_n814_ = \a[11]  ^ (((\a[14]  & ((new_n572_ & \a[17] ) | (~new_n572_ & ~\a[17] ) | ((~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))) & ((new_n572_ ^ \a[17] ) | (new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))) | ((~\a[14]  | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))) | ((~new_n572_ ^ \a[17] ) & (~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))) & (\a[14]  | ((new_n572_ ^ \a[17] ) ^ ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] ))))) & ((\a[14]  & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )) & (~new_n575_ | (new_n573_ ^ \a[17] ))) | (~new_n650_ & (~\a[14]  | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )) | (new_n575_ & (~new_n573_ ^ \a[17] ))) & (\a[14]  | (~new_n575_ ^ (new_n573_ ^ \a[17] ))))))) ^ (\a[14]  ^ (((new_n572_ & \a[17] ) | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] ))))) ^ (new_n571_ ^ \a[17] ))));
  assign new_n815_ = (new_n732_ ^ \a[11] ) ^ ((new_n733_ & \a[11] ) | ((~new_n733_ | ~\a[11] ) & (new_n733_ | \a[11] ) & (new_n734_ | (~new_n735_ & new_n806_))));
  assign new_n816_ = (new_n734_ | (~new_n735_ & new_n806_)) ^ (new_n733_ ^ \a[11] );
  assign new_n817_ = (~\a[8]  | (new_n735_ & ~new_n806_) | (~new_n735_ & new_n806_)) & ((\a[8]  & (~new_n735_ | new_n806_) & (new_n735_ | ~new_n806_)) | (~\a[8]  & (~new_n735_ ^ ~new_n806_)) | ((~new_n818_ | ~\a[8] ) & ((new_n818_ & \a[8] ) | (~new_n818_ & ~\a[8] ) | ((~new_n819_ | ~\a[8] ) & ((new_n819_ & \a[8] ) | (~new_n819_ & ~\a[8] ) | (~new_n820_ & (new_n821_ | ~new_n892_)))))));
  assign new_n818_ = (\a[11]  ^ (new_n655_ ^ ~new_n720_)) ^ ((new_n736_ & \a[11] ) | ((~new_n736_ | ~\a[11] ) & (new_n736_ | \a[11] ) & ((new_n737_ & \a[11] ) | ((~new_n737_ | ~\a[11] ) & (new_n737_ | \a[11] ) & (new_n738_ | (~new_n740_ & new_n805_))))));
  assign new_n819_ = (new_n736_ ^ \a[11] ) ^ ((new_n737_ & \a[11] ) | ((~new_n737_ | ~\a[11] ) & (new_n737_ | \a[11] ) & (new_n738_ | (~new_n740_ & new_n805_))));
  assign new_n820_ = \a[8]  & ((new_n737_ & \a[11] ) | (~new_n737_ & ~\a[11] ) | (~new_n738_ & (new_n740_ | ~new_n805_))) & ((new_n737_ ^ \a[11] ) | new_n738_ | (~new_n740_ & new_n805_));
  assign new_n821_ = (~\a[8]  | (new_n740_ & ~new_n805_) | (~new_n740_ & new_n805_)) & ((\a[8]  & (~new_n740_ | new_n805_) & (new_n740_ | ~new_n805_)) | (~\a[8]  & (~new_n740_ ^ ~new_n805_)) | ((~new_n822_ | ~\a[8] ) & ((new_n822_ & \a[8] ) | (~new_n822_ & ~\a[8] ) | ((~new_n823_ | ~\a[8] ) & ((new_n823_ & \a[8] ) | (~new_n823_ & ~\a[8] ) | (~new_n824_ & (new_n826_ | ~new_n891_)))))));
  assign new_n822_ = (new_n742_ ^ \a[11] ) ^ ((\a[11]  & ((new_n741_ & \a[14] ) | (~new_n741_ & ~\a[14] ) | ((new_n660_ | ~\a[14] ) & (((~new_n661_ | ~\a[14] ) & (new_n662_ | (new_n661_ & \a[14] ) | (~new_n661_ & ~\a[14] ))) | (~new_n660_ & \a[14] ) | (new_n660_ & ~\a[14] )))) & ((new_n741_ ^ \a[14] ) | (~new_n660_ & \a[14] ) | (((new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] ))) & (new_n660_ | ~\a[14] ) & (~new_n660_ | \a[14] )))) | (((\a[11]  & (((~new_n661_ | ~\a[14] ) & (new_n662_ | (new_n661_ & \a[14] ) | (~new_n661_ & ~\a[14] ))) | (~new_n660_ & \a[14] ) | (new_n660_ & ~\a[14] )) & ((new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] )) | (~new_n660_ ^ \a[14] ))) | (~new_n743_ & (~\a[11]  | (((new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] ))) & (new_n660_ | ~\a[14] ) & (~new_n660_ | \a[14] )) | ((~new_n661_ | ~\a[14] ) & (new_n662_ | (new_n661_ & \a[14] ) | (~new_n661_ & ~\a[14] )) & (new_n660_ ^ \a[14] ))) & (\a[11]  | (((new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] ))) ^ (~new_n660_ ^ \a[14] ))))) & (~\a[11]  | ((~new_n741_ | ~\a[14] ) & (new_n741_ | \a[14] ) & ((~new_n660_ & \a[14] ) | (((new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] ))) & (new_n660_ | ~\a[14] ) & (~new_n660_ | \a[14] )))) | ((~new_n741_ ^ \a[14] ) & (new_n660_ | ~\a[14] ) & (((~new_n661_ | ~\a[14] ) & (new_n662_ | (new_n661_ & \a[14] ) | (~new_n661_ & ~\a[14] ))) | (~new_n660_ & \a[14] ) | (new_n660_ & ~\a[14] )))) & (\a[11]  | ((new_n741_ ^ \a[14] ) ^ ((~new_n660_ & \a[14] ) | (((new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] ))) & (new_n660_ | ~\a[14] ) & (~new_n660_ | \a[14] )))))));
  assign new_n823_ = ((\a[11]  & ((~new_n660_ & \a[14] ) | (new_n660_ & ~\a[14] ) | ((~new_n661_ | ~\a[14] ) & (new_n662_ | (new_n661_ & \a[14] ) | (~new_n661_ & ~\a[14] )))) & ((~new_n660_ ^ \a[14] ) | (new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] )))) | (~new_n743_ & (~\a[11]  | ((new_n660_ | ~\a[14] ) & (~new_n660_ | \a[14] ) & ((new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] )))) | ((new_n660_ ^ \a[14] ) & (~new_n661_ | ~\a[14] ) & (new_n662_ | (new_n661_ & \a[14] ) | (~new_n661_ & ~\a[14] )))) & (\a[11]  | ((~new_n660_ ^ \a[14] ) ^ ((new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] ))))))) ^ (\a[11]  ^ ((~new_n741_ ^ ~\a[14] ) ^ ((~new_n660_ & \a[14] ) | ((new_n660_ | ~\a[14] ) & (~new_n660_ | \a[14] ) & ((new_n661_ & \a[14] ) | (~new_n662_ & (~new_n661_ | ~\a[14] ) & (new_n661_ | \a[14] )))))));
  assign new_n824_ = \a[8]  & (~new_n743_ | new_n825_) & (new_n743_ | ~new_n825_);
  assign new_n825_ = \a[11]  ^ ((~new_n660_ ^ \a[14] ) ^ ((new_n661_ & \a[14] ) | (~new_n662_ & (new_n661_ | \a[14] ) & (~new_n661_ | ~\a[14] ))));
  assign new_n826_ = (~new_n828_ | ~\a[8] ) & ((new_n828_ & \a[8] ) | (~new_n828_ & ~\a[8] ) | ((~\a[8]  | ((~new_n827_ | ~\a[11] ) & (new_n827_ | \a[11] ) & ((~new_n745_ & \a[11] ) | (((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] ))) & (new_n745_ | ~\a[11] ) & (~new_n745_ | \a[11] )))) | ((~new_n827_ ^ \a[11] ) & (new_n745_ | ~\a[11] ) & (((~new_n746_ | ~\a[11] ) & (new_n747_ | (new_n746_ & \a[11] ) | (~new_n746_ & ~\a[11] ))) | (~new_n745_ & \a[11] ) | (new_n745_ & ~\a[11] )))) & (((~\a[8]  | (((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] ))) & (new_n745_ | ~\a[11] ) & (~new_n745_ | \a[11] )) | ((~new_n746_ | ~\a[11] ) & (new_n747_ | (new_n746_ & \a[11] ) | (~new_n746_ & ~\a[11] )) & (new_n745_ ^ \a[11] ))) & (new_n829_ | (\a[8]  & (((~new_n746_ | ~\a[11] ) & (new_n747_ | (new_n746_ & \a[11] ) | (~new_n746_ & ~\a[11] ))) | (~new_n745_ & \a[11] ) | (new_n745_ & ~\a[11] )) & ((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] )) | (~new_n745_ ^ \a[11] ))) | (~\a[8]  & (((~new_n746_ | ~\a[11] ) & (new_n747_ | (new_n746_ & \a[11] ) | (~new_n746_ & ~\a[11] ))) ^ (~new_n745_ ^ \a[11] ))))) | (\a[8]  & ((new_n827_ & \a[11] ) | (~new_n827_ & ~\a[11] ) | ((new_n745_ | ~\a[11] ) & (((~new_n746_ | ~\a[11] ) & (new_n747_ | (new_n746_ & \a[11] ) | (~new_n746_ & ~\a[11] ))) | (~new_n745_ & \a[11] ) | (new_n745_ & ~\a[11] )))) & ((new_n827_ ^ \a[11] ) | (~new_n745_ & \a[11] ) | (((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] ))) & (new_n745_ | ~\a[11] ) & (~new_n745_ | \a[11] )))) | (~\a[8]  & ((~new_n827_ ^ \a[11] ) ^ ((~new_n745_ & \a[11] ) | (((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] ))) & (new_n745_ | ~\a[11] ) & (~new_n745_ | \a[11] ))))))));
  assign new_n827_ = ~new_n744_ ^ (new_n663_ ^ \a[14] );
  assign new_n828_ = (\a[11]  ^ ((new_n661_ ^ \a[14] ) ^ ((new_n663_ & \a[14] ) | (~new_n744_ & (~new_n663_ | ~\a[14] ) & (new_n663_ | \a[14] ))))) ^ ((\a[11]  & (new_n744_ | (new_n663_ & \a[14] ) | (~new_n663_ & ~\a[14] )) & (~new_n744_ | (new_n663_ ^ \a[14] ))) | ((~\a[11]  | (~new_n744_ & (~new_n663_ | ~\a[14] ) & (new_n663_ | \a[14] )) | (new_n744_ & (~new_n663_ ^ \a[14] ))) & (\a[11]  | (~new_n744_ ^ (new_n663_ ^ \a[14] ))) & ((~new_n745_ & \a[11] ) | ((new_n745_ | ~\a[11] ) & (~new_n745_ | \a[11] ) & ((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] )))))));
  assign new_n829_ = (~\a[8]  | ((~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] ) & ((new_n748_ & \a[11] ) | (~new_n830_ & (~new_n748_ | ~\a[11] ) & (new_n748_ | \a[11] )))) | ((~new_n746_ ^ \a[11] ) & (~new_n748_ | ~\a[11] ) & (new_n830_ | (new_n748_ & \a[11] ) | (~new_n748_ & ~\a[11] )))) & (((~\a[8]  | (~new_n830_ & (~new_n748_ | ~\a[11] ) & (new_n748_ | \a[11] )) | (new_n830_ & (~new_n748_ ^ \a[11] ))) & (((~new_n831_ | ~\a[8] ) & ((new_n831_ & \a[8] ) | (~new_n831_ & ~\a[8] ) | ((~new_n832_ | ~\a[8] ) & (new_n833_ | (new_n832_ & \a[8] ) | (~new_n832_ & ~\a[8] ))))) | (\a[8]  & (new_n830_ | (new_n748_ & \a[11] ) | (~new_n748_ & ~\a[11] )) & (~new_n830_ | (new_n748_ ^ \a[11] ))) | (~\a[8]  & (new_n830_ ^ (new_n748_ ^ \a[11] ))))) | (\a[8]  & ((new_n746_ & \a[11] ) | (~new_n746_ & ~\a[11] ) | ((~new_n748_ | ~\a[11] ) & (new_n830_ | (new_n748_ & \a[11] ) | (~new_n748_ & ~\a[11] )))) & ((new_n746_ ^ \a[11] ) | (new_n748_ & \a[11] ) | (~new_n830_ & (~new_n748_ | ~\a[11] ) & (new_n748_ | \a[11] )))) | (~\a[8]  & ((~new_n746_ ^ \a[11] ) ^ ((new_n748_ & \a[11] ) | (~new_n830_ & (~new_n748_ | ~\a[11] ) & (new_n748_ | \a[11] ))))));
  assign new_n830_ = ~new_n749_ & (new_n749_ | new_n803_ | ((new_n804_ | (~new_n674_ & new_n715_) | (new_n674_ & ~new_n715_)) & (new_n751_ | (~new_n804_ & (new_n674_ | ~new_n715_) & (~new_n674_ | new_n715_)) | (new_n804_ & (new_n674_ ^ new_n715_)))));
  assign new_n831_ = (~new_n749_ & ~new_n803_) ^ ((~new_n804_ & (new_n674_ | ~new_n715_) & (~new_n674_ | new_n715_)) | (~new_n751_ & (new_n804_ | (~new_n674_ & new_n715_) | (new_n674_ & ~new_n715_)) & (~new_n804_ | (~new_n674_ ^ new_n715_))));
  assign new_n832_ = ~new_n751_ ^ (~new_n804_ ^ (~new_n674_ ^ new_n715_));
  assign new_n833_ = (~new_n834_ | ~\a[8] ) & ((new_n834_ & \a[8] ) | (~new_n834_ & ~\a[8] ) | (~new_n835_ & (new_n835_ | new_n837_ | ((new_n890_ | (~new_n759_ & new_n800_) | (new_n759_ & ~new_n800_)) & (new_n838_ | (~new_n890_ & (new_n759_ | ~new_n800_) & (~new_n759_ | new_n800_)) | (new_n890_ & (new_n759_ ^ new_n800_)))))));
  assign new_n834_ = (new_n752_ ^ ~new_n802_) ^ (new_n754_ | (new_n801_ & (new_n756_ | (~new_n759_ & new_n800_))));
  assign new_n835_ = ~new_n836_ & (~new_n801_ | (~new_n756_ & (new_n759_ | ~new_n800_))) & (new_n801_ | new_n756_ | (~new_n759_ & new_n800_));
  assign new_n836_ = \a[8]  ^ (~\b[19]  | (((\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (new_n201_ | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ))));
  assign new_n837_ = new_n836_ & (~new_n801_ ^ (new_n756_ | (~new_n759_ & new_n800_)));
  assign new_n838_ = (~new_n839_ | new_n889_) & ((new_n839_ & ~new_n889_) | (~new_n839_ & new_n889_) | (~new_n841_ & (~new_n888_ | (~new_n843_ & (new_n846_ | ~new_n887_)))));
  assign new_n839_ = new_n840_ ^ (new_n761_ | (((~new_n799_ & (new_n686_ | ~new_n709_) & (~new_n686_ | new_n709_)) | (~new_n763_ & (new_n799_ | (~new_n686_ & new_n709_) | (new_n686_ & ~new_n709_)) & (~new_n799_ | (~new_n686_ ^ new_n709_)))) & ~new_n761_ & ~new_n797_));
  assign new_n840_ = ~new_n798_ ^ ((new_n681_ | (new_n710_ & (new_n683_ | (~new_n686_ & new_n709_)))) ^ (new_n679_ ^ ~new_n711_));
  assign new_n841_ = ~new_n842_ & (new_n761_ | new_n797_ | ((new_n799_ | (~new_n686_ & new_n709_) | (new_n686_ & ~new_n709_)) & (new_n763_ | (~new_n799_ & (new_n686_ | ~new_n709_) & (~new_n686_ | new_n709_)) | (new_n799_ & (new_n686_ ^ new_n709_))))) & ((~new_n761_ & ~new_n797_) | (~new_n799_ & (new_n686_ | ~new_n709_) & (~new_n686_ | new_n709_)) | (~new_n763_ & (new_n799_ | (~new_n686_ & new_n709_) | (new_n686_ & ~new_n709_)) & (~new_n799_ | (~new_n686_ ^ new_n709_))));
  assign new_n842_ = \a[8]  ^ ((~new_n199_ | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[17]  | (\a[5]  ^ \a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[18]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[16]  | (\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n843_ = ~new_n845_ & (~new_n763_ | new_n844_) & (new_n763_ | ~new_n844_);
  assign new_n844_ = ~new_n799_ ^ (new_n686_ ^ ~new_n709_);
  assign new_n845_ = \a[8]  ^ ((~new_n144_ | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[16]  | (\a[5]  ^ \a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[17]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[15]  | (\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n846_ = (~new_n847_ | new_n885_) & ((new_n847_ & ~new_n885_) | (~new_n847_ & new_n885_) | (~new_n848_ & (new_n848_ | new_n884_ | ((new_n886_ | (~new_n771_ & new_n794_) | (new_n771_ & ~new_n794_)) & (new_n850_ | (~new_n886_ & (new_n771_ | ~new_n794_) & (~new_n771_ | new_n794_)) | (new_n886_ & (new_n771_ ^ new_n794_)))))));
  assign new_n847_ = (new_n764_ ^ ~new_n796_) ^ (new_n766_ | (new_n795_ & (new_n768_ | (~new_n771_ & new_n794_))));
  assign new_n848_ = ~new_n849_ & (~new_n795_ | (~new_n768_ & (new_n771_ | ~new_n794_))) & (new_n795_ | new_n768_ | (~new_n771_ & new_n794_));
  assign new_n849_ = \a[8]  ^ ((((~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] ) & ((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )))) | ((~\b[14]  ^ \b[15] ) & (~\b[13]  | ~\b[14] ) & (new_n142_ | (\b[13]  & \b[14] ) | (~\b[13]  & ~\b[14] ))) | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[14]  | (\a[5]  ^ \a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[15]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[13]  | (\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n850_ = (~new_n851_ | new_n883_) & ((new_n851_ & ~new_n883_) | (~new_n851_ & new_n883_) | (~new_n853_ & (~new_n882_ | (~new_n855_ & (new_n858_ | ~new_n881_)))));
  assign new_n851_ = new_n852_ ^ (new_n774_ | (new_n790_ & ((~new_n793_ & (new_n697_ | (~new_n696_ & new_n704_) | (new_n696_ & ~new_n704_)) & (~new_n697_ | (~new_n696_ ^ new_n704_))) | (~new_n776_ & (new_n793_ | (~new_n697_ & (new_n696_ | ~new_n704_) & (~new_n696_ | new_n704_)) | (new_n697_ & (new_n696_ ^ new_n704_))) & (~new_n793_ | (~new_n697_ ^ (~new_n696_ ^ new_n704_)))))));
  assign new_n852_ = ~new_n791_ ^ ((new_n692_ ^ ~new_n693_) ^ ((new_n694_ & ~new_n695_) | ((~new_n694_ | new_n695_) & (new_n694_ | ~new_n695_) & ((~new_n696_ & new_n704_) | (~new_n697_ & (new_n696_ | ~new_n704_) & (~new_n696_ | new_n704_))))));
  assign new_n853_ = ~new_n854_ & (~new_n790_ | ((new_n793_ | (~new_n697_ & (new_n696_ | ~new_n704_) & (~new_n696_ | new_n704_)) | (new_n697_ & (new_n696_ ^ new_n704_))) & (new_n776_ | (~new_n793_ & (new_n697_ | (~new_n696_ & new_n704_) | (new_n696_ & ~new_n704_)) & (~new_n697_ | (~new_n696_ ^ new_n704_))) | (new_n793_ & (new_n697_ ^ (~new_n696_ ^ new_n704_)))))) & (new_n790_ | (~new_n793_ & (new_n697_ | (~new_n696_ & new_n704_) | (new_n696_ & ~new_n704_)) & (~new_n697_ | (~new_n696_ ^ new_n704_))) | (~new_n776_ & (new_n793_ | (~new_n697_ & (new_n696_ | ~new_n704_) & (~new_n696_ | new_n704_)) | (new_n697_ & (new_n696_ ^ new_n704_))) & (~new_n793_ | (~new_n697_ ^ (~new_n696_ ^ new_n704_)))));
  assign new_n854_ = \a[8]  ^ ((~new_n107_ | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[11]  | (\a[5]  ^ \a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[12]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[10]  | (\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n855_ = ~new_n857_ & (~new_n776_ | new_n856_) & (new_n776_ | ~new_n856_);
  assign new_n856_ = ~new_n793_ ^ (~new_n697_ ^ (~new_n696_ ^ new_n704_));
  assign new_n857_ = \a[8]  ^ ((~new_n135_ | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[10]  | (\a[5]  ^ \a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[11]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[9]  | (\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n858_ = (~new_n860_ | new_n878_) & ((~new_n861_ & (~new_n877_ | ((new_n880_ | (new_n859_ & ~new_n782_) | (~new_n859_ & new_n782_)) & (new_n863_ | (~new_n880_ & (~new_n859_ | new_n782_) & (new_n859_ | ~new_n782_)) | (new_n880_ & (~new_n859_ ^ ~new_n782_)))))) | (new_n860_ & ~new_n878_) | (~new_n860_ & new_n878_));
  assign new_n859_ = new_n781_ ^ ~new_n789_;
  assign new_n860_ = (new_n777_ ^ ~new_n778_) ^ ((new_n779_ & ~new_n780_) | (((~new_n781_ & new_n789_) | (~new_n782_ & (new_n781_ | ~new_n789_) & (~new_n781_ | new_n789_))) & (~new_n779_ | new_n780_) & (new_n779_ | ~new_n780_)));
  assign new_n861_ = ~new_n862_ & ((new_n779_ & ~new_n780_) | (~new_n779_ & new_n780_) | ((new_n781_ | ~new_n789_) & (new_n782_ | (~new_n781_ & new_n789_) | (new_n781_ & ~new_n789_)))) & ((new_n779_ ^ ~new_n780_) | (~new_n781_ & new_n789_) | (~new_n782_ & (new_n781_ | ~new_n789_) & (~new_n781_ | new_n789_)));
  assign new_n862_ = \a[8]  ^ ((((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))) | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[8]  | (\a[5]  ^ \a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[9]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[7]  | (\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n863_ = (~new_n864_ | new_n865_) & ((new_n864_ & ~new_n865_) | (~new_n864_ & new_n865_) | ((~new_n866_ | new_n867_) & (((new_n868_ | ~new_n876_) & (new_n869_ | (~new_n868_ & new_n876_) | (new_n868_ & ~new_n876_))) | (new_n866_ & ~new_n867_) | (~new_n866_ & new_n867_))));
  assign new_n864_ = (new_n786_ | (~new_n787_ & new_n788_)) ^ (new_n785_ ^ (~\a[11]  ^ (new_n784_ & (~new_n98_ | ~new_n783_))));
  assign new_n865_ = \a[8]  ^ ((~new_n88_ | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[6]  | (\a[5]  ^ \a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[7]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[5]  | (\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n866_ = new_n787_ ^ ~new_n788_;
  assign new_n867_ = \a[8]  ^ ((~new_n91_ | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[5]  | (\a[5]  ^ \a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[6]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[4]  | (\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n868_ = \a[8]  ^ ((~new_n94_ | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[4]  | (\a[5]  ^ \a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[5]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[3]  | (\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n869_ = (~new_n872_ | (\a[8]  ^ (new_n871_ & (~new_n98_ | ~new_n870_)))) & ((~new_n873_ & (new_n874_ | ~new_n875_)) | (new_n872_ & (~\a[8]  ^ (new_n871_ & (~new_n98_ | ~new_n870_)))) | (~new_n872_ & (~\a[8]  | ~new_n871_ | (new_n98_ & new_n870_)) & (\a[8]  | (new_n871_ & (~new_n98_ | ~new_n870_)))));
  assign new_n870_ = (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (~\a[7]  | ~\a[8] ) & (\a[7]  | \a[8] );
  assign new_n871_ = (~\b[3]  | (~\a[5]  ^ ~\a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[4]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[2]  | (\a[6]  ^ \a[7] ) | (~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ));
  assign new_n872_ = ((\b[0]  & (\a[8]  ^ ~\a[9] ) & (~\a[9]  | ~\a[10] ) & (\a[9]  | \a[10] )) | (\b[1]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (~\a[10]  ^ \a[11] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (~\a[10]  | ~\a[11] ) & (\a[10]  | \a[11] ))) ^ (\a[11]  & \b[0]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ));
  assign new_n873_ = \b[0]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] ) & (~\b[0]  | (~\a[5]  ^ ~\a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[1]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  ^ \a[8] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[0]  | (\a[6]  ^ \a[7] ) | (~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[1]  | (~\a[5]  ^ ~\a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[2]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  ^ \a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )));
  assign new_n874_ = \a[8]  ^ (((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (~\a[5]  ^ ~\a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[3]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[1]  | (\a[6]  ^ \a[7] ) | (~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n875_ = (\b[0]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] )) ^ ((~\b[0]  | (~\a[5]  ^ ~\a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[1]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  ^ \a[8] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[0]  | (\a[6]  ^ \a[7] ) | (~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[1]  | (~\a[5]  ^ ~\a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[2]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  ^ \a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n876_ = (~\a[11]  | ((~\b[0]  | (~\a[8]  ^ ~\a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[1]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  ^ \a[11] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )))) ^ ((~\b[1]  | (~\a[8]  ^ ~\a[9] ) | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] )) & (~\b[2]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  ^ \a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (\a[9]  ^ \a[10] ) | (~\a[8]  ^ ~\a[9] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] )));
  assign new_n877_ = ~new_n862_ ^ ((new_n779_ ^ ~new_n780_) ^ ((~new_n781_ & new_n789_) | (~new_n782_ & (new_n781_ | ~new_n789_) & (~new_n781_ | new_n789_))));
  assign new_n878_ = \a[8]  ^ (new_n879_ & (~new_n870_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n879_ = (~\b[9]  | (~\a[5]  ^ ~\a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[10]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[8]  | (\a[6]  ^ \a[7] ) | (~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ));
  assign new_n880_ = \a[8]  ^ ((~\b[7]  | (\a[5]  ^ \a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[8]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[6]  | (\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & ((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n79_ & (~\b[7]  ^ \b[8] ))));
  assign new_n881_ = ~new_n857_ ^ (new_n776_ ^ ~new_n856_);
  assign new_n882_ = ~new_n854_ ^ (new_n790_ ^ ((~new_n793_ & (new_n697_ | (~new_n696_ & new_n704_) | (new_n696_ & ~new_n704_)) & (~new_n697_ | (~new_n696_ ^ new_n704_))) | (~new_n776_ & (new_n793_ | (~new_n697_ & (new_n696_ | ~new_n704_) & (~new_n696_ | new_n704_)) | (new_n697_ & (new_n696_ ^ new_n704_))) & (~new_n793_ | (~new_n697_ ^ (~new_n696_ ^ new_n704_))))));
  assign new_n883_ = \a[8]  ^ ((~new_n133_ | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[12]  | (\a[5]  ^ \a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[13]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[11]  | (\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n884_ = new_n849_ & (~new_n795_ ^ (new_n768_ | (~new_n771_ & new_n794_)));
  assign new_n885_ = \a[8]  ^ ((~new_n186_ | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[15]  | (\a[5]  ^ \a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[16]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[14]  | (\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n886_ = \a[8]  ^ ((~\b[13]  | (\a[5]  ^ \a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[14]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[12]  | (\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & ((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n142_ & (~\b[13]  ^ \b[14] ))));
  assign new_n887_ = ~new_n845_ ^ (new_n763_ ^ ~new_n844_);
  assign new_n888_ = ~new_n842_ ^ ((~new_n761_ & ~new_n797_) ^ ((~new_n799_ & (new_n686_ | ~new_n709_) & (~new_n686_ | new_n709_)) | (~new_n763_ & (new_n799_ | (~new_n686_ & new_n709_) | (new_n686_ & ~new_n709_)) & (~new_n799_ | (~new_n686_ ^ new_n709_)))));
  assign new_n889_ = \a[8]  ^ ((~new_n253_ | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & (~\b[18]  | (\a[5]  ^ \a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[19]  | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  ^ \a[8] )) & (~\b[17]  | (\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n890_ = \a[8]  ^ (((\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~new_n201_ ^ ~\b[19] )) & (~\b[19]  | (\a[5]  ^ \a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[18]  | (\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n891_ = \a[8]  ^ (new_n743_ ^ ~new_n825_);
  assign new_n892_ = \a[8]  ^ ((new_n737_ ^ \a[11] ) ^ (new_n738_ | (~new_n740_ & new_n805_)));
  assign new_n893_ = (~new_n649_ ^ ~\a[14] ) ^ ((\a[14]  & ((new_n571_ & \a[17] ) | (~new_n571_ & ~\a[17] ) | ((~new_n572_ | ~\a[17] ) & ((new_n572_ & \a[17] ) | (~new_n572_ & ~\a[17] ) | ((~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))))) & ((new_n571_ ^ \a[17] ) | (new_n572_ & \a[17] ) | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))))) | ((~\a[14]  | ((~new_n571_ | ~\a[17] ) & (new_n571_ | \a[17] ) & ((new_n572_ & \a[17] ) | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))))) | ((~new_n571_ ^ \a[17] ) & (~new_n572_ | ~\a[17] ) & ((new_n572_ & \a[17] ) | (~new_n572_ & ~\a[17] ) | ((~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))))) & (\a[14]  | ((new_n571_ ^ \a[17] ) ^ ((new_n572_ & \a[17] ) | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] ))))))) & ((\a[14]  & ((new_n572_ & \a[17] ) | (~new_n572_ & ~\a[17] ) | ((~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))) & ((new_n572_ ^ \a[17] ) | (new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))) | ((~\a[14]  | ((~new_n572_ | ~\a[17] ) & (new_n572_ | \a[17] ) & ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )))) | ((~new_n572_ ^ \a[17] ) & (~new_n573_ | ~\a[17] ) & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )))) & (\a[14]  | ((new_n572_ ^ \a[17] ) ^ ((new_n573_ & \a[17] ) | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] ))))) & ((\a[14]  & (new_n575_ | (new_n573_ & \a[17] ) | (~new_n573_ & ~\a[17] )) & (~new_n575_ | (new_n573_ ^ \a[17] ))) | (~new_n650_ & (~\a[14]  | (~new_n575_ & (~new_n573_ | ~\a[17] ) & (new_n573_ | \a[17] )) | (new_n575_ & (~new_n573_ ^ \a[17] ))) & (\a[14]  | (~new_n575_ ^ (new_n573_ ^ \a[17] )))))))));
  assign new_n894_ = (new_n896_ ^ \a[14] ) ^ ((\a[14]  & ((new_n895_ & \a[17] ) | (~new_n895_ & ~\a[17] ) | ((~new_n562_ | ~\a[17] ) & ((new_n562_ & \a[17] ) | (~new_n562_ & ~\a[17] ) | ((~new_n563_ | ~\a[17] ) & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )))))) & ((new_n895_ ^ \a[17] ) | (new_n562_ & \a[17] ) | ((~new_n562_ | ~\a[17] ) & (new_n562_ | \a[17] ) & ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )))))) | ((~\a[14]  | ((~new_n895_ | ~\a[17] ) & (new_n895_ | \a[17] ) & ((new_n562_ & \a[17] ) | ((~new_n562_ | ~\a[17] ) & (new_n562_ | \a[17] ) & ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )))))) | ((~new_n895_ ^ \a[17] ) & (~new_n562_ | ~\a[17] ) & ((new_n562_ & \a[17] ) | (~new_n562_ & ~\a[17] ) | ((~new_n563_ | ~\a[17] ) & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )))))) & (\a[14]  | ((new_n895_ ^ \a[17] ) ^ ((new_n562_ & \a[17] ) | ((~new_n562_ | ~\a[17] ) & (new_n562_ | \a[17] ) & ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] ))))))) & ((\a[14]  & ((new_n562_ & \a[17] ) | (~new_n562_ & ~\a[17] ) | ((~new_n563_ | ~\a[17] ) & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )))) & ((new_n562_ ^ \a[17] ) | (new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )))) | ((~\a[14]  | ((~new_n562_ | ~\a[17] ) & (new_n562_ | \a[17] ) & ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )))) | ((~new_n562_ ^ \a[17] ) & (~new_n563_ | ~\a[17] ) & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )))) & (\a[14]  | ((new_n562_ ^ \a[17] ) ^ ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] ))))) & ((\a[14]  & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )) & (~new_n564_ | (new_n563_ ^ \a[17] ))) | (~new_n643_ & (~\a[14]  | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )) | (new_n564_ & (~new_n563_ ^ \a[17] ))) & (\a[14]  | (~new_n564_ ^ (new_n563_ ^ \a[17] )))))))));
  assign new_n895_ = ~new_n68_ ^ (new_n531_ ^ \a[20] );
  assign new_n896_ = (\a[17]  ^ ((~new_n560_ ^ \a[20] ) ^ ((~new_n531_ | ~\a[20] ) & (new_n68_ | (new_n531_ & \a[20] ) | (~new_n531_ & ~\a[20] ))))) ^ ((\a[17]  & (new_n68_ | (new_n531_ & \a[20] ) | (~new_n531_ & ~\a[20] )) & (~new_n68_ | (new_n531_ ^ \a[20] ))) | ((~\a[17]  | (~new_n68_ & (~new_n531_ | ~\a[20] ) & (new_n531_ | \a[20] )) | (new_n68_ & (~new_n531_ ^ \a[20] ))) & (\a[17]  | (~new_n68_ ^ (new_n531_ ^ \a[20] ))) & ((new_n562_ & \a[17] ) | ((new_n562_ | \a[17] ) & (~new_n562_ | ~\a[17] ) & ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )))))));
  assign new_n897_ = ((\a[14]  & ((new_n562_ & \a[17] ) | (~new_n562_ & ~\a[17] ) | ((~new_n563_ | ~\a[17] ) & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )))) & ((new_n562_ ^ \a[17] ) | (new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )))) | (((\a[14]  & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )) & (~new_n564_ | (new_n563_ ^ \a[17] ))) | (~new_n643_ & (~\a[14]  | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )) | (new_n564_ & (~new_n563_ ^ \a[17] ))) & (\a[14]  | (~new_n564_ ^ (new_n563_ ^ \a[17] ))))) & (~\a[14]  | ((~new_n562_ | ~\a[17] ) & (new_n562_ | \a[17] ) & ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )))) | ((~new_n562_ ^ \a[17] ) & (~new_n563_ | ~\a[17] ) & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )))) & (\a[14]  | ((new_n562_ ^ \a[17] ) ^ ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] ))))))) ^ (\a[14]  ^ ((~new_n895_ ^ ~\a[17] ) ^ ((new_n562_ & \a[17] ) | ((~new_n562_ | ~\a[17] ) & (new_n562_ | \a[17] ) & ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )))))));
  assign new_n898_ = (~\a[11]  | (new_n722_ & ((new_n642_ & \a[14] ) | (~new_n643_ & (~new_n642_ | ~\a[14] ) & (new_n642_ | \a[14] )))) | (~new_n722_ & (~new_n642_ | ~\a[14] ) & (new_n643_ | (new_n642_ & \a[14] ) | (~new_n642_ & ~\a[14] )))) & (((~\a[11]  | (~new_n643_ & (~new_n642_ | ~\a[14] ) & (new_n642_ | \a[14] )) | (new_n643_ & (~new_n642_ ^ \a[14] ))) & (((~new_n723_ | ~\a[11] ) & (((~new_n724_ | ~\a[11] ) & (new_n725_ | (~new_n724_ & ~\a[11] ) | (new_n724_ & \a[11] ))) | (new_n723_ & \a[11] ) | (~new_n723_ & ~\a[11] ))) | (\a[11]  & (new_n643_ | (new_n642_ & \a[14] ) | (~new_n642_ & ~\a[14] )) & (~new_n643_ | (new_n642_ ^ \a[14] ))) | (~\a[11]  & (new_n643_ ^ (new_n642_ ^ \a[14] ))))) | (\a[11]  & (~new_n722_ | ((~new_n642_ | ~\a[14] ) & (new_n643_ | (new_n642_ & \a[14] ) | (~new_n642_ & ~\a[14] )))) & (new_n722_ | (new_n642_ & \a[14] ) | (~new_n643_ & (~new_n642_ | ~\a[14] ) & (new_n642_ | \a[14] )))) | (~\a[11]  & (~new_n722_ ^ ((new_n642_ & \a[14] ) | (~new_n643_ & (~new_n642_ | ~\a[14] ) & (new_n642_ | \a[14] ))))));
  assign new_n899_ = (~new_n896_ | ~\a[14] ) & ((new_n896_ & \a[14] ) | (~new_n896_ & ~\a[14] ) | ((~\a[14]  | ((~new_n895_ | ~\a[17] ) & (new_n895_ | \a[17] ) & ((new_n562_ & \a[17] ) | ((~new_n562_ | ~\a[17] ) & (new_n562_ | \a[17] ) & ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )))))) | ((~new_n895_ ^ \a[17] ) & (~new_n562_ | ~\a[17] ) & ((new_n562_ & \a[17] ) | (~new_n562_ & ~\a[17] ) | ((~new_n563_ | ~\a[17] ) & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )))))) & ((\a[14]  & ((new_n895_ & \a[17] ) | (~new_n895_ & ~\a[17] ) | ((~new_n562_ | ~\a[17] ) & ((new_n562_ & \a[17] ) | (~new_n562_ & ~\a[17] ) | ((~new_n563_ | ~\a[17] ) & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )))))) & ((new_n895_ ^ \a[17] ) | (new_n562_ & \a[17] ) | ((~new_n562_ | ~\a[17] ) & (new_n562_ | \a[17] ) & ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )))))) | (~\a[14]  & ((~new_n895_ ^ \a[17] ) ^ ((new_n562_ & \a[17] ) | ((~new_n562_ | ~\a[17] ) & (new_n562_ | \a[17] ) & ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] ))))))) | ((~\a[14]  | ((~new_n562_ | ~\a[17] ) & (new_n562_ | \a[17] ) & ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )))) | ((~new_n562_ ^ \a[17] ) & (~new_n563_ | ~\a[17] ) & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )))) & ((\a[14]  & ((new_n562_ & \a[17] ) | (~new_n562_ & ~\a[17] ) | ((~new_n563_ | ~\a[17] ) & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )))) & ((new_n562_ ^ \a[17] ) | (new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )))) | (~\a[14]  & ((~new_n562_ ^ \a[17] ) ^ ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] ))))) | ((~\a[14]  | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )) | (new_n564_ & (~new_n563_ ^ \a[17] ))) & (new_n643_ | (\a[14]  & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )) & (~new_n564_ | (new_n563_ ^ \a[17] ))) | (~\a[14]  & (new_n564_ ^ (new_n563_ ^ \a[17] ))))))))));
  assign new_n900_ = (new_n901_ ^ new_n902_) ^ (~new_n904_ ^ ((~\a[14]  | (~new_n66_ & new_n561_) | (new_n66_ & ~new_n561_)) & (new_n899_ | (\a[14]  & (new_n66_ | ~new_n561_) & (~new_n66_ | new_n561_)) | (~\a[14]  & (new_n66_ ^ new_n561_)))));
  assign new_n901_ = \a[23]  ^ ((new_n546_ & \a[26] ) | ((new_n546_ | \a[26] ) & (~new_n546_ | ~\a[26] ) & ((new_n557_ & \a[26] ) | ((~new_n557_ | ~\a[26] ) & (new_n557_ | \a[26] ) & ((new_n532_ & \a[26] ) | ((~new_n532_ | ~\a[26] ) & (new_n532_ | \a[26] ) & ((new_n521_ & \a[26] ) | (~new_n520_ & (new_n521_ | \a[26] ) & (~new_n521_ | ~\a[26] )))))))));
  assign new_n902_ = (~new_n903_ ^ ~\a[26] ) ^ ((~new_n552_ | ~\a[32] ) & ((new_n552_ & \a[32] ) | (~new_n552_ & ~\a[32] ) | (~new_n547_ & (~new_n556_ | ((~new_n535_ | ~\a[32] ) & (new_n534_ | (new_n535_ & \a[32] ) | (~new_n535_ & ~\a[32] )))))));
  assign new_n903_ = (~\a[29]  | ((~new_n552_ | ~\a[32] ) & (new_n552_ | \a[32] ) & (new_n547_ | (new_n556_ & ((new_n535_ & \a[32] ) | (~new_n534_ & (~new_n535_ | ~\a[32] ) & (new_n535_ | \a[32] )))))) | ((~new_n552_ ^ \a[32] ) & ~new_n547_ & (~new_n556_ | ((~new_n535_ | ~\a[32] ) & (new_n534_ | (new_n535_ & \a[32] ) | (~new_n535_ & ~\a[32] )))))) & (((~\a[29]  | (new_n556_ & ((new_n535_ & \a[32] ) | (~new_n534_ & (~new_n535_ | ~\a[32] ) & (new_n535_ | \a[32] )))) | (~new_n556_ & (~new_n535_ | ~\a[32] ) & (new_n534_ | (new_n535_ & \a[32] ) | (~new_n535_ & ~\a[32] )))) & (((~\a[29]  | (~new_n534_ & (~new_n535_ | ~\a[32] ) & (new_n535_ | \a[32] )) | (new_n534_ & (~new_n535_ ^ \a[32] ))) & (new_n533_ | (\a[29]  & (new_n534_ | (new_n535_ & \a[32] ) | (~new_n535_ & ~\a[32] )) & (~new_n534_ | (new_n535_ ^ \a[32] ))) | (~\a[29]  & (new_n534_ ^ (new_n535_ ^ \a[32] ))))) | (\a[29]  & (~new_n556_ | ((~new_n535_ | ~\a[32] ) & (new_n534_ | (new_n535_ & \a[32] ) | (~new_n535_ & ~\a[32] )))) & (new_n556_ | (new_n535_ & \a[32] ) | (~new_n534_ & (~new_n535_ | ~\a[32] ) & (new_n535_ | \a[32] )))) | (~\a[29]  & (~new_n556_ ^ ((new_n535_ & \a[32] ) | (~new_n534_ & (~new_n535_ | ~\a[32] ) & (new_n535_ | \a[32] ))))))) | (\a[29]  & ((new_n552_ & \a[32] ) | (~new_n552_ & ~\a[32] ) | (~new_n547_ & (~new_n556_ | ((~new_n535_ | ~\a[32] ) & (new_n534_ | (new_n535_ & \a[32] ) | (~new_n535_ & ~\a[32] )))))) & ((new_n552_ ^ \a[32] ) | new_n547_ | (new_n556_ & ((new_n535_ & \a[32] ) | (~new_n534_ & (~new_n535_ | ~\a[32] ) & (new_n535_ | \a[32] )))))) | (~\a[29]  & ((~new_n552_ ^ \a[32] ) ^ (new_n547_ | (new_n556_ & ((new_n535_ & \a[32] ) | (~new_n534_ & (~new_n535_ | ~\a[32] ) & (new_n535_ | \a[32] ))))))));
  assign new_n904_ = (new_n553_ | ((\a[38]  & ~\b[18] ) ^ (~\b[19]  | (((\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (\a[36]  ^ \a[37] ) | (\a[35]  ^ \a[36] )) & (new_n201_ | (\a[37]  & \a[38] ) | (~\a[37]  & ~\a[38] ) | (\a[35]  & \a[36] ) | (~\a[35]  & ~\a[36] )))))) & (~\a[38]  | ~\b[18]  | (\b[19]  & (((~\a[37]  | ~\a[38] ) & (\a[37]  | \a[38] ) & (~\a[36]  ^ \a[37] ) & (~\a[35]  ^ \a[36] )) | (~new_n201_ & (~\a[37]  | ~\a[38] ) & (\a[37]  | \a[38] ) & (~\a[35]  | ~\a[36] ) & (\a[35]  | \a[36] )))));
  assign new_n905_ = (\a[38]  & ~\b[19] ) ^ (((new_n545_ & \a[23] ) | ((~new_n545_ | ~\a[23] ) & (new_n545_ | \a[23] ) & ((new_n559_ & \a[23] ) | (~new_n558_ & (~new_n559_ | ~\a[23] ) & (new_n559_ | \a[23] ))))) ^ (\a[20]  ^ ~\a[35] ));
  assign new_n906_ = ~new_n1006_ ^ (\a[2]  ^ ((new_n907_ & \a[5] ) | (~new_n908_ & (~new_n907_ | ~\a[5] ) & (new_n907_ | \a[5] ))));
  assign new_n907_ = ((\a[8]  & ((new_n894_ & \a[11] ) | (~new_n894_ & ~\a[11] ) | ((~new_n897_ | ~\a[11] ) & (new_n898_ | (new_n897_ & \a[11] ) | (~new_n897_ & ~\a[11] )))) & ((new_n894_ ^ \a[11] ) | (new_n897_ & \a[11] ) | (~new_n898_ & (~new_n897_ | ~\a[11] ) & (new_n897_ | \a[11] )))) | ((~\a[8]  | ((~new_n894_ | ~\a[11] ) & (new_n894_ | \a[11] ) & ((new_n897_ & \a[11] ) | (~new_n898_ & (~new_n897_ | ~\a[11] ) & (new_n897_ | \a[11] )))) | ((~new_n894_ ^ \a[11] ) & (~new_n897_ | ~\a[11] ) & (new_n898_ | (new_n897_ & \a[11] ) | (~new_n897_ & ~\a[11] )))) & (\a[8]  | ((new_n894_ ^ \a[11] ) ^ ((new_n897_ & \a[11] ) | (~new_n898_ & (~new_n897_ | ~\a[11] ) & (new_n897_ | \a[11] ))))) & ((\a[8]  & (new_n898_ | (new_n897_ & \a[11] ) | (~new_n897_ & ~\a[11] )) & (~new_n898_ | (new_n897_ ^ \a[11] ))) | (~new_n640_ & (~\a[8]  | (~new_n898_ & (~new_n897_ | ~\a[11] ) & (new_n897_ | \a[11] )) | (new_n898_ & (~new_n897_ ^ \a[11] ))) & (\a[8]  | (~new_n898_ ^ (new_n897_ ^ \a[11] ))))))) ^ (\a[8]  ^ (((new_n894_ & \a[11] ) | ((~new_n894_ | ~\a[11] ) & (new_n894_ | \a[11] ) & ((new_n897_ & \a[11] ) | (~new_n898_ & (~new_n897_ | ~\a[11] ) & (new_n897_ | \a[11] ))))) ^ (\a[11]  ^ (new_n65_ ^ ~new_n899_))));
  assign new_n908_ = (~\a[5]  | (new_n912_ & (new_n909_ | (~new_n640_ & new_n911_))) | (~new_n912_ & ~new_n909_ & (new_n640_ | ~new_n911_))) & (((~\a[5]  | (~new_n640_ & new_n911_) | (new_n640_ & ~new_n911_)) & (((~new_n913_ | ~\a[5] ) & ((new_n913_ & \a[5] ) | (~new_n913_ & ~\a[5] ) | ((~new_n914_ | ~\a[5] ) & (new_n915_ | (new_n914_ & \a[5] ) | (~new_n914_ & ~\a[5] ))))) | (\a[5]  & (new_n640_ | ~new_n911_) & (~new_n640_ | new_n911_)) | (~\a[5]  & (new_n640_ ^ new_n911_)))) | (\a[5]  & (~new_n912_ | (~new_n909_ & (new_n640_ | ~new_n911_))) & (new_n912_ | new_n909_ | (~new_n640_ & new_n911_))) | (~\a[5]  & (~new_n912_ ^ (new_n909_ | (~new_n640_ & new_n911_)))));
  assign new_n909_ = \a[8]  & (~new_n898_ | new_n910_) & (new_n898_ | ~new_n910_);
  assign new_n910_ = \a[11]  ^ (((\a[14]  & ((new_n562_ & \a[17] ) | (~new_n562_ & ~\a[17] ) | ((~new_n563_ | ~\a[17] ) & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )))) & ((new_n562_ ^ \a[17] ) | (new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )))) | ((~\a[14]  | ((~new_n562_ | ~\a[17] ) & (new_n562_ | \a[17] ) & ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )))) | ((~new_n562_ ^ \a[17] ) & (~new_n563_ | ~\a[17] ) & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )))) & (\a[14]  | ((new_n562_ ^ \a[17] ) ^ ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] ))))) & ((\a[14]  & (new_n564_ | (new_n563_ & \a[17] ) | (~new_n563_ & ~\a[17] )) & (~new_n564_ | (new_n563_ ^ \a[17] ))) | (~new_n643_ & (~\a[14]  | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] )) | (new_n564_ & (~new_n563_ ^ \a[17] ))) & (\a[14]  | (~new_n564_ ^ (new_n563_ ^ \a[17] ))))))) ^ (\a[14]  ^ (((new_n562_ & \a[17] ) | ((~new_n562_ | ~\a[17] ) & (new_n562_ | \a[17] ) & ((new_n563_ & \a[17] ) | (~new_n564_ & (~new_n563_ | ~\a[17] ) & (new_n563_ | \a[17] ))))) ^ (new_n895_ ^ \a[17] ))));
  assign new_n911_ = \a[8]  ^ (new_n898_ ^ ~new_n910_);
  assign new_n912_ = \a[8]  ^ ((new_n894_ ^ \a[11] ) ^ ((new_n897_ & \a[11] ) | (~new_n898_ & (new_n897_ | \a[11] ) & (~new_n897_ | ~\a[11] ))));
  assign new_n913_ = ((\a[8]  & ((new_n641_ & \a[11] ) | (~new_n641_ & ~\a[11] ) | ((~new_n723_ | ~\a[11] ) & ((new_n723_ & \a[11] ) | (~new_n723_ & ~\a[11] ) | ((~new_n724_ | ~\a[11] ) & (new_n725_ | (new_n724_ & \a[11] ) | (~new_n724_ & ~\a[11] )))))) & ((new_n641_ ^ \a[11] ) | (new_n723_ & \a[11] ) | ((~new_n723_ | ~\a[11] ) & (new_n723_ | \a[11] ) & ((new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] )))))) | (((\a[8]  & ((new_n723_ & \a[11] ) | (~new_n723_ & ~\a[11] ) | ((~new_n724_ | ~\a[11] ) & (new_n725_ | (new_n724_ & \a[11] ) | (~new_n724_ & ~\a[11] )))) & ((new_n723_ ^ \a[11] ) | (new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] )))) | ((~\a[8]  | ((~new_n723_ | ~\a[11] ) & (new_n723_ | \a[11] ) & ((new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] )))) | ((~new_n723_ ^ \a[11] ) & (~new_n724_ | ~\a[11] ) & (new_n725_ | (new_n724_ & \a[11] ) | (~new_n724_ & ~\a[11] )))) & (\a[8]  | ((new_n723_ ^ \a[11] ) ^ ((new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] ))))) & ((\a[8]  & (new_n725_ | (new_n724_ & \a[11] ) | (~new_n724_ & ~\a[11] )) & (~new_n725_ | (new_n724_ ^ \a[11] ))) | (~new_n807_ & (~\a[8]  | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] )) | (new_n725_ & (~new_n724_ ^ \a[11] ))) & (\a[8]  | (~new_n725_ ^ (new_n724_ ^ \a[11] ))))))) & (~\a[8]  | ((~new_n641_ | ~\a[11] ) & (new_n641_ | \a[11] ) & ((new_n723_ & \a[11] ) | ((~new_n723_ | ~\a[11] ) & (new_n723_ | \a[11] ) & ((new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] )))))) | ((~new_n641_ ^ \a[11] ) & (~new_n723_ | ~\a[11] ) & ((new_n723_ & \a[11] ) | (~new_n723_ & ~\a[11] ) | ((~new_n724_ | ~\a[11] ) & (new_n725_ | (new_n724_ & \a[11] ) | (~new_n724_ & ~\a[11] )))))) & (\a[8]  | ((new_n641_ ^ \a[11] ) ^ ((new_n723_ & \a[11] ) | ((~new_n723_ | ~\a[11] ) & (new_n723_ | \a[11] ) & ((new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] ))))))))) ^ (new_n721_ ^ \a[8] );
  assign new_n914_ = ((\a[8]  & ((new_n723_ & \a[11] ) | (~new_n723_ & ~\a[11] ) | ((~new_n724_ | ~\a[11] ) & (new_n725_ | (new_n724_ & \a[11] ) | (~new_n724_ & ~\a[11] )))) & ((new_n723_ ^ \a[11] ) | (new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] )))) | (((\a[8]  & (new_n725_ | (new_n724_ & \a[11] ) | (~new_n724_ & ~\a[11] )) & (~new_n725_ | (new_n724_ ^ \a[11] ))) | (~new_n807_ & (~\a[8]  | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] )) | (new_n725_ & (~new_n724_ ^ \a[11] ))) & (\a[8]  | (~new_n725_ ^ (new_n724_ ^ \a[11] ))))) & (~\a[8]  | ((~new_n723_ | ~\a[11] ) & (new_n723_ | \a[11] ) & ((new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] )))) | ((~new_n723_ ^ \a[11] ) & (~new_n724_ | ~\a[11] ) & (new_n725_ | (new_n724_ & \a[11] ) | (~new_n724_ & ~\a[11] )))) & (\a[8]  | ((new_n723_ ^ \a[11] ) ^ ((new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] ))))))) ^ (\a[8]  ^ ((~new_n641_ ^ ~\a[11] ) ^ ((new_n723_ & \a[11] ) | ((~new_n723_ | ~\a[11] ) & (new_n723_ | \a[11] ) & ((new_n724_ & \a[11] ) | (~new_n725_ & (~new_n724_ | ~\a[11] ) & (new_n724_ | \a[11] )))))));
  assign new_n915_ = (~\a[5]  | (new_n918_ & (new_n916_ | (~new_n807_ & new_n917_))) | (~new_n918_ & ~new_n916_ & (new_n807_ | ~new_n917_))) & (((~\a[5]  | (~new_n807_ & new_n917_) | (new_n807_ & ~new_n917_)) & (((~new_n919_ | ~\a[5] ) & ((new_n919_ & \a[5] ) | (~new_n919_ & ~\a[5] ) | ((~new_n920_ | ~\a[5] ) & (new_n921_ | (new_n920_ & \a[5] ) | (~new_n920_ & ~\a[5] ))))) | (\a[5]  & (new_n807_ | ~new_n917_) & (~new_n807_ | new_n917_)) | (~\a[5]  & (new_n807_ ^ new_n917_)))) | (\a[5]  & (~new_n918_ | (~new_n916_ & (new_n807_ | ~new_n917_))) & (new_n918_ | new_n916_ | (~new_n807_ & new_n917_))) | (~\a[5]  & (~new_n918_ ^ (new_n916_ | (~new_n807_ & new_n917_)))));
  assign new_n916_ = \a[8]  & (new_n725_ | (~new_n724_ & ~\a[11] ) | (new_n724_ & \a[11] )) & (~new_n725_ | (~new_n724_ ^ ~\a[11] ));
  assign new_n917_ = \a[8]  ^ (~new_n725_ ^ (~new_n724_ ^ ~\a[11] ));
  assign new_n918_ = \a[8]  ^ ((new_n723_ ^ \a[11] ) ^ ((new_n724_ & \a[11] ) | (~new_n725_ & (new_n724_ | \a[11] ) & (~new_n724_ | ~\a[11] ))));
  assign new_n919_ = (~new_n808_ ^ ~\a[8] ) ^ ((new_n809_ & \a[8] ) | ((~new_n809_ | ~\a[8] ) & (new_n809_ | \a[8] ) & ((\a[8]  & ((new_n893_ & \a[11] ) | (~new_n893_ & ~\a[11] ) | ((~new_n727_ | ~\a[11] ) & (new_n728_ | (new_n727_ & \a[11] ) | (~new_n727_ & ~\a[11] )))) & ((new_n893_ ^ \a[11] ) | (new_n727_ & \a[11] ) | (~new_n728_ & (~new_n727_ | ~\a[11] ) & (new_n727_ | \a[11] )))) | (~new_n810_ & (~\a[8]  | ((~new_n893_ | ~\a[11] ) & (new_n893_ | \a[11] ) & ((new_n727_ & \a[11] ) | (~new_n728_ & (~new_n727_ | ~\a[11] ) & (new_n727_ | \a[11] )))) | ((~new_n893_ ^ \a[11] ) & (~new_n727_ | ~\a[11] ) & (new_n728_ | (new_n727_ & \a[11] ) | (~new_n727_ & ~\a[11] )))) & (\a[8]  | ((new_n893_ ^ \a[11] ) ^ ((new_n727_ & \a[11] ) | (~new_n728_ & (~new_n727_ | ~\a[11] ) & (new_n727_ | \a[11] )))))))));
  assign new_n920_ = (~new_n809_ ^ ~\a[8] ) ^ ((\a[8]  & ((new_n893_ & \a[11] ) | (~new_n893_ & ~\a[11] ) | ((~new_n727_ | ~\a[11] ) & (new_n728_ | ~new_n814_))) & ((new_n893_ ^ \a[11] ) | (new_n727_ & \a[11] ) | (~new_n728_ & new_n814_))) | (~new_n810_ & (~\a[8]  | ((~new_n893_ | ~\a[11] ) & (new_n893_ | \a[11] ) & ((new_n727_ & \a[11] ) | (~new_n728_ & new_n814_))) | ((~new_n893_ ^ \a[11] ) & (~new_n727_ | ~\a[11] ) & (new_n728_ | ~new_n814_))) & (\a[8]  | ((new_n893_ ^ \a[11] ) ^ ((new_n727_ & \a[11] ) | (~new_n728_ & new_n814_))))));
  assign new_n921_ = (~\a[5]  | (new_n810_ & ~new_n922_) | (~new_n810_ & new_n922_)) & (((~new_n923_ | ~\a[5] ) & ((new_n923_ & \a[5] ) | (~new_n923_ & ~\a[5] ) | ((~new_n924_ | ~\a[5] ) & (((~new_n925_ | ~\a[5] ) & (new_n926_ | (~new_n925_ & ~\a[5] ) | (new_n925_ & \a[5] ))) | (new_n924_ & \a[5] ) | (~new_n924_ & ~\a[5] ))))) | (\a[5]  & (~new_n810_ | new_n922_) & (new_n810_ | ~new_n922_)) | (~\a[5]  & (~new_n810_ ^ ~new_n922_)));
  assign new_n922_ = \a[8]  ^ ((new_n893_ ^ \a[11] ) ^ ((new_n727_ & \a[11] ) | (~new_n728_ & (new_n727_ | \a[11] ) & (~new_n727_ | ~\a[11] ))));
  assign new_n923_ = ((\a[8]  & (new_n812_ | ~new_n813_) & (~new_n812_ | new_n813_)) | (((new_n815_ & \a[8] ) | ((~new_n815_ | ~\a[8] ) & (new_n815_ | \a[8] ) & ((new_n816_ & \a[8] ) | (~new_n817_ & (~new_n816_ | ~\a[8] ) & (new_n816_ | \a[8] ))))) & (~\a[8]  | (~new_n812_ & new_n813_) | (new_n812_ & ~new_n813_)) & (\a[8]  | (~new_n812_ ^ new_n813_)))) ^ (\a[8]  ^ (new_n814_ ^ (new_n811_ | (~new_n812_ & new_n813_))));
  assign new_n924_ = ((new_n815_ & \a[8] ) | ((new_n815_ | \a[8] ) & (~new_n815_ | ~\a[8] ) & ((new_n816_ & \a[8] ) | (~new_n817_ & (~new_n816_ | ~\a[8] ) & (new_n816_ | \a[8] ))))) ^ (\a[8]  ^ (new_n812_ ^ ~new_n813_));
  assign new_n925_ = (~new_n815_ ^ ~\a[8] ) ^ ((new_n816_ & \a[8] ) | (~new_n817_ & (new_n816_ | \a[8] ) & (~new_n816_ | ~\a[8] )));
  assign new_n926_ = (~\a[5]  | (~new_n817_ & (~new_n816_ | ~\a[8] ) & (new_n816_ | \a[8] )) | (new_n817_ & (~new_n816_ ^ \a[8] ))) & (((~new_n927_ | ~\a[5] ) & ((new_n927_ & \a[5] ) | (~new_n927_ & ~\a[5] ) | ((~new_n928_ | ~\a[5] ) & (((~new_n929_ | ~\a[5] ) & (new_n930_ | (~new_n929_ & ~\a[5] ) | (new_n929_ & \a[5] ))) | (new_n928_ & \a[5] ) | (~new_n928_ & ~\a[5] ))))) | (\a[5]  & (new_n817_ | (new_n816_ & \a[8] ) | (~new_n816_ & ~\a[8] )) & (~new_n817_ | (new_n816_ ^ \a[8] ))) | (~\a[5]  & (new_n817_ ^ (new_n816_ ^ \a[8] ))));
  assign new_n927_ = (\a[8]  ^ (new_n735_ ^ ~new_n806_)) ^ ((new_n818_ & \a[8] ) | ((~new_n818_ | ~\a[8] ) & (new_n818_ | \a[8] ) & ((new_n819_ & \a[8] ) | ((~new_n819_ | ~\a[8] ) & (new_n819_ | \a[8] ) & (new_n820_ | (~new_n821_ & new_n892_))))));
  assign new_n928_ = (new_n818_ ^ \a[8] ) ^ ((new_n819_ & \a[8] ) | ((~new_n819_ | ~\a[8] ) & (new_n819_ | \a[8] ) & (new_n820_ | (~new_n821_ & new_n892_))));
  assign new_n929_ = (new_n820_ | (~new_n821_ & new_n892_)) ^ (new_n819_ ^ \a[8] );
  assign new_n930_ = (~\a[5]  | (new_n821_ & ~new_n892_) | (~new_n821_ & new_n892_)) & ((\a[5]  & (~new_n821_ | new_n892_) & (new_n821_ | ~new_n892_)) | (~\a[5]  & (~new_n821_ ^ ~new_n892_)) | ((~new_n931_ | ~\a[5] ) & ((new_n931_ & \a[5] ) | (~new_n931_ & ~\a[5] ) | ((~new_n932_ | ~\a[5] ) & ((new_n932_ & \a[5] ) | (~new_n932_ & ~\a[5] ) | (~new_n933_ & (new_n934_ | ~new_n1005_)))))));
  assign new_n931_ = (\a[8]  ^ (new_n740_ ^ ~new_n805_)) ^ ((new_n822_ & \a[8] ) | ((~new_n822_ | ~\a[8] ) & (new_n822_ | \a[8] ) & ((new_n823_ & \a[8] ) | ((~new_n823_ | ~\a[8] ) & (new_n823_ | \a[8] ) & (new_n824_ | (~new_n826_ & new_n891_))))));
  assign new_n932_ = (new_n822_ ^ \a[8] ) ^ ((new_n823_ & \a[8] ) | ((~new_n823_ | ~\a[8] ) & (new_n823_ | \a[8] ) & (new_n824_ | (~new_n826_ & new_n891_))));
  assign new_n933_ = \a[5]  & ((new_n823_ & \a[8] ) | (~new_n823_ & ~\a[8] ) | (~new_n824_ & (new_n826_ | ~new_n891_))) & ((new_n823_ ^ \a[8] ) | new_n824_ | (~new_n826_ & new_n891_));
  assign new_n934_ = (~\a[5]  | (new_n826_ & ~new_n891_) | (~new_n826_ & new_n891_)) & ((\a[5]  & (~new_n826_ | new_n891_) & (new_n826_ | ~new_n891_)) | (~\a[5]  & (~new_n826_ ^ ~new_n891_)) | ((~new_n935_ | ~\a[5] ) & ((new_n935_ & \a[5] ) | (~new_n935_ & ~\a[5] ) | ((~new_n936_ | ~\a[5] ) & ((new_n936_ & \a[5] ) | (~new_n936_ & ~\a[5] ) | ((~\a[5]  | (~new_n829_ & new_n1004_) | (new_n829_ & ~new_n1004_)) & (new_n937_ | (\a[5]  & (new_n829_ | ~new_n1004_) & (~new_n829_ | new_n1004_)) | (~\a[5]  & (new_n829_ ^ new_n1004_)))))))));
  assign new_n935_ = (new_n828_ ^ \a[8] ) ^ ((\a[8]  & ((new_n827_ & \a[11] ) | (~new_n827_ & ~\a[11] ) | ((new_n745_ | ~\a[11] ) & (((~new_n746_ | ~\a[11] ) & (new_n747_ | (new_n746_ & \a[11] ) | (~new_n746_ & ~\a[11] ))) | (~new_n745_ & \a[11] ) | (new_n745_ & ~\a[11] )))) & ((new_n827_ ^ \a[11] ) | (~new_n745_ & \a[11] ) | (((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] ))) & (new_n745_ | ~\a[11] ) & (~new_n745_ | \a[11] )))) | (((\a[8]  & (((~new_n746_ | ~\a[11] ) & (new_n747_ | (new_n746_ & \a[11] ) | (~new_n746_ & ~\a[11] ))) | (~new_n745_ & \a[11] ) | (new_n745_ & ~\a[11] )) & ((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] )) | (~new_n745_ ^ \a[11] ))) | (~new_n829_ & (~\a[8]  | (((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] ))) & (new_n745_ | ~\a[11] ) & (~new_n745_ | \a[11] )) | ((~new_n746_ | ~\a[11] ) & (new_n747_ | (new_n746_ & \a[11] ) | (~new_n746_ & ~\a[11] )) & (new_n745_ ^ \a[11] ))) & (\a[8]  | (((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] ))) ^ (~new_n745_ ^ \a[11] ))))) & (~\a[8]  | ((~new_n827_ | ~\a[11] ) & (new_n827_ | \a[11] ) & ((~new_n745_ & \a[11] ) | (((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] ))) & (new_n745_ | ~\a[11] ) & (~new_n745_ | \a[11] )))) | ((~new_n827_ ^ \a[11] ) & (new_n745_ | ~\a[11] ) & (((~new_n746_ | ~\a[11] ) & (new_n747_ | (new_n746_ & \a[11] ) | (~new_n746_ & ~\a[11] ))) | (~new_n745_ & \a[11] ) | (new_n745_ & ~\a[11] )))) & (\a[8]  | ((new_n827_ ^ \a[11] ) ^ ((~new_n745_ & \a[11] ) | (((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] ))) & (new_n745_ | ~\a[11] ) & (~new_n745_ | \a[11] )))))));
  assign new_n936_ = ((\a[8]  & ((~new_n745_ & \a[11] ) | (new_n745_ & ~\a[11] ) | ((~new_n746_ | ~\a[11] ) & (new_n747_ | (new_n746_ & \a[11] ) | (~new_n746_ & ~\a[11] )))) & ((~new_n745_ ^ \a[11] ) | (new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] )))) | (~new_n829_ & (~\a[8]  | ((new_n745_ | ~\a[11] ) & (~new_n745_ | \a[11] ) & ((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] )))) | ((new_n745_ ^ \a[11] ) & (~new_n746_ | ~\a[11] ) & (new_n747_ | (new_n746_ & \a[11] ) | (~new_n746_ & ~\a[11] )))) & (\a[8]  | ((~new_n745_ ^ \a[11] ) ^ ((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] ))))))) ^ (\a[8]  ^ ((~new_n827_ ^ ~\a[11] ) ^ ((~new_n745_ & \a[11] ) | ((new_n745_ | ~\a[11] ) & (~new_n745_ | \a[11] ) & ((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] )))))));
  assign new_n937_ = (~new_n939_ | ~\a[5] ) & ((new_n939_ & \a[5] ) | (~new_n939_ & ~\a[5] ) | ((~\a[5]  | ((~new_n938_ | ~\a[8] ) & (new_n938_ | \a[8] ) & ((new_n831_ & \a[8] ) | ((~new_n831_ | ~\a[8] ) & (new_n831_ | \a[8] ) & ((new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] )))))) | ((~new_n938_ ^ \a[8] ) & (~new_n831_ | ~\a[8] ) & ((new_n831_ & \a[8] ) | (~new_n831_ & ~\a[8] ) | ((~new_n832_ | ~\a[8] ) & (new_n833_ | (new_n832_ & \a[8] ) | (~new_n832_ & ~\a[8] )))))) & ((\a[5]  & ((new_n938_ & \a[8] ) | (~new_n938_ & ~\a[8] ) | ((~new_n831_ | ~\a[8] ) & ((new_n831_ & \a[8] ) | (~new_n831_ & ~\a[8] ) | ((~new_n832_ | ~\a[8] ) & (new_n833_ | (new_n832_ & \a[8] ) | (~new_n832_ & ~\a[8] )))))) & ((new_n938_ ^ \a[8] ) | (new_n831_ & \a[8] ) | ((~new_n831_ | ~\a[8] ) & (new_n831_ | \a[8] ) & ((new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] )))))) | (~\a[5]  & ((~new_n938_ ^ \a[8] ) ^ ((new_n831_ & \a[8] ) | ((~new_n831_ | ~\a[8] ) & (new_n831_ | \a[8] ) & ((new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] ))))))) | ((~\a[5]  | ((~new_n831_ | ~\a[8] ) & (new_n831_ | \a[8] ) & ((new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] )))) | ((~new_n831_ ^ \a[8] ) & (~new_n832_ | ~\a[8] ) & (new_n833_ | (new_n832_ & \a[8] ) | (~new_n832_ & ~\a[8] )))) & (new_n940_ | (\a[5]  & ((new_n831_ & \a[8] ) | (~new_n831_ & ~\a[8] ) | ((~new_n832_ | ~\a[8] ) & (new_n833_ | (new_n832_ & \a[8] ) | (~new_n832_ & ~\a[8] )))) & ((new_n831_ ^ \a[8] ) | (new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] )))) | (~\a[5]  & ((~new_n831_ ^ \a[8] ) ^ ((new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] ))))))))));
  assign new_n938_ = ~new_n830_ ^ (new_n748_ ^ \a[11] );
  assign new_n939_ = ((\a[8]  & (new_n830_ | (new_n748_ & \a[11] ) | (~new_n748_ & ~\a[11] )) & (~new_n830_ | (new_n748_ ^ \a[11] ))) | (((new_n831_ & \a[8] ) | ((~new_n831_ | ~\a[8] ) & (new_n831_ | \a[8] ) & ((new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] ))))) & (~\a[8]  | (~new_n830_ & (~new_n748_ | ~\a[11] ) & (new_n748_ | \a[11] )) | (new_n830_ & (~new_n748_ ^ \a[11] ))) & (\a[8]  | (~new_n830_ ^ (new_n748_ ^ \a[11] ))))) ^ (\a[8]  ^ ((new_n746_ ^ \a[11] ) ^ ((new_n748_ & \a[11] ) | (~new_n830_ & (~new_n748_ | ~\a[11] ) & (new_n748_ | \a[11] )))));
  assign new_n940_ = (~\a[5]  | ((~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] ) & ((new_n834_ & \a[8] ) | (~new_n941_ & (~new_n834_ | ~\a[8] ) & (new_n834_ | \a[8] )))) | ((~new_n832_ ^ \a[8] ) & (~new_n834_ | ~\a[8] ) & (new_n941_ | (new_n834_ & \a[8] ) | (~new_n834_ & ~\a[8] )))) & (((~\a[5]  | (~new_n941_ & (~new_n834_ | ~\a[8] ) & (new_n834_ | \a[8] )) | (new_n941_ & (~new_n834_ ^ \a[8] ))) & (((~new_n942_ | ~\a[5] ) & ((new_n942_ & \a[5] ) | (~new_n942_ & ~\a[5] ) | ((~new_n943_ | ~\a[5] ) & (new_n945_ | (new_n943_ & \a[5] ) | (~new_n943_ & ~\a[5] ))))) | (\a[5]  & (new_n941_ | (new_n834_ & \a[8] ) | (~new_n834_ & ~\a[8] )) & (~new_n941_ | (new_n834_ ^ \a[8] ))) | (~\a[5]  & (new_n941_ ^ (new_n834_ ^ \a[8] ))))) | (\a[5]  & ((new_n832_ & \a[8] ) | (~new_n832_ & ~\a[8] ) | ((~new_n834_ | ~\a[8] ) & (new_n941_ | (new_n834_ & \a[8] ) | (~new_n834_ & ~\a[8] )))) & ((new_n832_ ^ \a[8] ) | (new_n834_ & \a[8] ) | (~new_n941_ & (~new_n834_ | ~\a[8] ) & (new_n834_ | \a[8] )))) | (~\a[5]  & ((~new_n832_ ^ \a[8] ) ^ ((new_n834_ & \a[8] ) | (~new_n941_ & (~new_n834_ | ~\a[8] ) & (new_n834_ | \a[8] ))))));
  assign new_n941_ = ~new_n835_ & (new_n835_ | new_n837_ | ((new_n890_ | (~new_n759_ & new_n800_) | (new_n759_ & ~new_n800_)) & (new_n838_ | (~new_n890_ & (new_n759_ | ~new_n800_) & (~new_n759_ | new_n800_)) | (new_n890_ & (new_n759_ ^ new_n800_)))));
  assign new_n942_ = (~new_n835_ & ~new_n837_) ^ ((~new_n890_ & (new_n759_ | ~new_n800_) & (~new_n759_ | new_n800_)) | (~new_n838_ & (new_n890_ | (~new_n759_ & new_n800_) | (new_n759_ & ~new_n800_)) & (~new_n890_ | (~new_n759_ ^ new_n800_))));
  assign new_n943_ = new_n838_ ^ ~new_n944_;
  assign new_n944_ = ~new_n890_ ^ (new_n759_ ^ ~new_n800_);
  assign new_n945_ = (~new_n946_ | ~\a[5] ) & ((new_n946_ & \a[5] ) | (~new_n946_ & ~\a[5] ) | (~new_n947_ & (new_n947_ | new_n1002_ | ((new_n1003_ | (~new_n846_ & new_n887_) | (new_n846_ & ~new_n887_)) & (new_n949_ | (~new_n1003_ & (new_n846_ | ~new_n887_) & (~new_n846_ | new_n887_)) | (new_n1003_ & (new_n846_ ^ new_n887_)))))));
  assign new_n946_ = (new_n839_ ^ ~new_n889_) ^ (new_n841_ | (new_n888_ & (new_n843_ | (~new_n846_ & new_n887_))));
  assign new_n947_ = ~new_n948_ & (~new_n888_ | (~new_n843_ & (new_n846_ | ~new_n887_))) & (new_n888_ | new_n843_ | (~new_n846_ & new_n887_));
  assign new_n948_ = \a[5]  ^ (~\b[19]  | (((\a[3]  ^ \a[4] ) | (\a[2]  ^ \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (new_n201_ | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ))));
  assign new_n949_ = (~new_n950_ | new_n1001_) & ((new_n950_ & ~new_n1001_) | (~new_n950_ & new_n1001_) | (~new_n952_ & (~new_n1000_ | (~new_n954_ & (new_n957_ | ~new_n999_)))));
  assign new_n950_ = new_n951_ ^ (new_n848_ | (((~new_n886_ & (new_n771_ | ~new_n794_) & (~new_n771_ | new_n794_)) | (~new_n850_ & (new_n886_ | (~new_n771_ & new_n794_) | (new_n771_ & ~new_n794_)) & (~new_n886_ | (~new_n771_ ^ new_n794_)))) & ~new_n848_ & ~new_n884_));
  assign new_n951_ = ~new_n885_ ^ ((new_n766_ | (new_n795_ & (new_n768_ | (~new_n771_ & new_n794_)))) ^ (new_n764_ ^ ~new_n796_));
  assign new_n952_ = ~new_n953_ & (new_n848_ | new_n884_ | ((new_n886_ | (~new_n771_ & new_n794_) | (new_n771_ & ~new_n794_)) & (new_n850_ | (~new_n886_ & (new_n771_ | ~new_n794_) & (~new_n771_ | new_n794_)) | (new_n886_ & (new_n771_ ^ new_n794_))))) & ((~new_n848_ & ~new_n884_) | (~new_n886_ & (new_n771_ | ~new_n794_) & (~new_n771_ | new_n794_)) | (~new_n850_ & (new_n886_ | (~new_n771_ & new_n794_) | (new_n771_ & ~new_n794_)) & (~new_n886_ | (~new_n771_ ^ new_n794_))));
  assign new_n953_ = \a[5]  ^ ((~new_n199_ | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[17]  | (\a[2]  ^ \a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[18]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[16]  | (\a[3]  ^ \a[4] ) | (\a[2]  ^ \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n954_ = ~new_n956_ & (~new_n850_ | new_n955_) & (new_n850_ | ~new_n955_);
  assign new_n955_ = ~new_n886_ ^ (new_n771_ ^ ~new_n794_);
  assign new_n956_ = \a[5]  ^ ((~new_n144_ | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[16]  | (\a[2]  ^ \a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[17]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[15]  | (\a[3]  ^ \a[4] ) | (\a[2]  ^ \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n957_ = (~new_n958_ | new_n997_) & ((new_n958_ & ~new_n997_) | (~new_n958_ & new_n997_) | (~new_n959_ & (new_n959_ | new_n996_ | ((new_n998_ | (~new_n858_ & new_n881_) | (new_n858_ & ~new_n881_)) & (new_n961_ | (~new_n998_ & (new_n858_ | ~new_n881_) & (~new_n858_ | new_n881_)) | (new_n998_ & (new_n858_ ^ new_n881_)))))));
  assign new_n958_ = (new_n851_ ^ ~new_n883_) ^ (new_n853_ | (new_n882_ & (new_n855_ | (~new_n858_ & new_n881_))));
  assign new_n959_ = ~new_n960_ & (~new_n882_ | (~new_n855_ & (new_n858_ | ~new_n881_))) & (new_n882_ | new_n855_ | (~new_n858_ & new_n881_));
  assign new_n960_ = \a[5]  ^ ((((~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] ) & ((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )))) | ((~\b[14]  ^ \b[15] ) & (~\b[13]  | ~\b[14] ) & (new_n142_ | (\b[13]  & \b[14] ) | (~\b[13]  & ~\b[14] ))) | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[14]  | (\a[2]  ^ \a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[15]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[13]  | (\a[3]  ^ \a[4] ) | (\a[2]  ^ \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n961_ = (~new_n962_ | new_n995_) & ((new_n962_ & ~new_n995_) | (~new_n962_ & new_n995_) | (~new_n964_ & (~new_n994_ | (~new_n966_ & (new_n969_ | ~new_n993_)))));
  assign new_n962_ = new_n963_ ^ (new_n861_ | (new_n877_ & ((~new_n880_ & (new_n782_ | (~new_n781_ & new_n789_) | (new_n781_ & ~new_n789_)) & (~new_n782_ | (~new_n781_ ^ new_n789_))) | (~new_n863_ & (new_n880_ | (~new_n782_ & (new_n781_ | ~new_n789_) & (~new_n781_ | new_n789_)) | (new_n782_ & (new_n781_ ^ new_n789_))) & (~new_n880_ | (~new_n782_ ^ (~new_n781_ ^ new_n789_)))))));
  assign new_n963_ = ~new_n878_ ^ ((new_n777_ ^ ~new_n778_) ^ ((new_n779_ & ~new_n780_) | ((~new_n779_ | new_n780_) & (new_n779_ | ~new_n780_) & ((~new_n781_ & new_n789_) | (~new_n782_ & (new_n781_ | ~new_n789_) & (~new_n781_ | new_n789_))))));
  assign new_n964_ = ~new_n965_ & (~new_n877_ | ((new_n880_ | (~new_n782_ & (new_n781_ | ~new_n789_) & (~new_n781_ | new_n789_)) | (new_n782_ & (new_n781_ ^ new_n789_))) & (new_n863_ | (~new_n880_ & (new_n782_ | (~new_n781_ & new_n789_) | (new_n781_ & ~new_n789_)) & (~new_n782_ | (~new_n781_ ^ new_n789_))) | (new_n880_ & (new_n782_ ^ (~new_n781_ ^ new_n789_)))))) & (new_n877_ | (~new_n880_ & (new_n782_ | (~new_n781_ & new_n789_) | (new_n781_ & ~new_n789_)) & (~new_n782_ | (~new_n781_ ^ new_n789_))) | (~new_n863_ & (new_n880_ | (~new_n782_ & (new_n781_ | ~new_n789_) & (~new_n781_ | new_n789_)) | (new_n782_ & (new_n781_ ^ new_n789_))) & (~new_n880_ | (~new_n782_ ^ (~new_n781_ ^ new_n789_)))));
  assign new_n965_ = \a[5]  ^ ((~new_n107_ | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[11]  | (\a[2]  ^ \a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[12]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[10]  | (\a[3]  ^ \a[4] ) | (\a[2]  ^ \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n966_ = ~new_n968_ & (~new_n863_ | new_n967_) & (new_n863_ | ~new_n967_);
  assign new_n967_ = ~new_n880_ ^ (~new_n782_ ^ (~new_n781_ ^ new_n789_));
  assign new_n968_ = \a[5]  ^ ((~new_n135_ | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[10]  | (\a[2]  ^ \a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[11]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[9]  | (\a[3]  ^ \a[4] ) | (\a[2]  ^ \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n969_ = (~new_n971_ | new_n990_) & ((new_n971_ & ~new_n990_) | (~new_n971_ & new_n990_) | (~new_n972_ & (~new_n974_ | ((new_n992_ | (new_n970_ & ~new_n869_) | (~new_n970_ & new_n869_)) & (new_n975_ | (~new_n992_ & (~new_n970_ | new_n869_) & (new_n970_ | ~new_n869_)) | (new_n992_ & (~new_n970_ ^ ~new_n869_)))))));
  assign new_n970_ = new_n868_ ^ ~new_n876_;
  assign new_n971_ = (new_n864_ ^ ~new_n865_) ^ ((new_n866_ & ~new_n867_) | (((~new_n868_ & new_n876_) | (~new_n869_ & (new_n868_ | ~new_n876_) & (~new_n868_ | new_n876_))) & (~new_n866_ | new_n867_) & (new_n866_ | ~new_n867_)));
  assign new_n972_ = ~new_n973_ & ((new_n866_ & ~new_n867_) | (~new_n866_ & new_n867_) | ((new_n868_ | ~new_n876_) & (new_n869_ | (~new_n868_ & new_n876_) | (new_n868_ & ~new_n876_)))) & ((new_n866_ ^ ~new_n867_) | (~new_n868_ & new_n876_) | (~new_n869_ & (new_n868_ | ~new_n876_) & (~new_n868_ | new_n876_)));
  assign new_n973_ = \a[5]  ^ ((((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))) | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[8]  | (\a[2]  ^ \a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[9]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[7]  | (\a[3]  ^ \a[4] ) | (\a[2]  ^ \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n974_ = ~new_n973_ ^ ((new_n866_ ^ ~new_n867_) ^ ((~new_n868_ & new_n876_) | (~new_n869_ & (new_n868_ | ~new_n876_) & (~new_n868_ | new_n876_))));
  assign new_n975_ = (~new_n976_ | new_n977_) & ((new_n976_ & ~new_n977_) | (~new_n976_ & new_n977_) | ((~new_n978_ | new_n979_) & (((new_n980_ | ~new_n989_) & (new_n983_ | (~new_n980_ & new_n989_) | (new_n980_ & ~new_n989_))) | (new_n978_ & ~new_n979_) | (~new_n978_ & new_n979_))));
  assign new_n976_ = (new_n873_ | (~new_n874_ & new_n875_)) ^ (new_n872_ ^ (~\a[8]  ^ (new_n871_ & (~new_n98_ | ~new_n870_))));
  assign new_n977_ = \a[5]  ^ ((~new_n88_ | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[6]  | (\a[2]  ^ \a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[7]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[5]  | (\a[3]  ^ \a[4] ) | (\a[2]  ^ \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n978_ = new_n874_ ^ ~new_n875_;
  assign new_n979_ = \a[5]  ^ ((~new_n91_ | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[5]  | (\a[2]  ^ \a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[6]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[4]  | (\a[3]  ^ \a[4] ) | (\a[2]  ^ \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n980_ = \a[5]  ^ (new_n982_ & (~new_n94_ | ~new_n981_));
  assign new_n981_ = (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (~\a[4]  | ~\a[5] ) & (\a[4]  | \a[5] );
  assign new_n982_ = (~\b[4]  | (~\a[2]  ^ ~\a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[5]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[3]  | (\a[3]  ^ \a[4] ) | (~\a[2]  ^ ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ));
  assign new_n983_ = (~new_n985_ | (\a[5]  ^ (new_n984_ & (~new_n98_ | ~new_n981_)))) & ((~new_n986_ & (new_n987_ | ~new_n988_)) | (new_n985_ & (~\a[5]  ^ (new_n984_ & (~new_n98_ | ~new_n981_)))) | (~new_n985_ & (~\a[5]  | ~new_n984_ | (new_n98_ & new_n981_)) & (\a[5]  | (new_n984_ & (~new_n98_ | ~new_n981_)))));
  assign new_n984_ = (~\b[3]  | (~\a[2]  ^ ~\a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[4]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[2]  | (\a[3]  ^ \a[4] ) | (~\a[2]  ^ ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ));
  assign new_n985_ = ((\b[0]  & (\a[5]  ^ ~\a[6] ) & (~\a[6]  | ~\a[7] ) & (\a[6]  | \a[7] )) | (\b[1]  & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (~\a[7]  ^ \a[8] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (~\a[7]  | ~\a[8] ) & (\a[7]  | \a[8] ))) ^ (\a[8]  & \b[0]  & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ));
  assign new_n986_ = \b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (~\b[0]  | (~\a[2]  ^ ~\a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[1]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  ^ \a[5] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[0]  | (\a[3]  ^ \a[4] ) | (~\a[2]  ^ ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[1]  | (~\a[2]  ^ ~\a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[2]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  ^ \a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )));
  assign new_n987_ = \a[5]  ^ (((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (~\a[2]  ^ ~\a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[3]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[1]  | (\a[3]  ^ \a[4] ) | (~\a[2]  ^ ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n988_ = (\b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] )) ^ ((~\b[0]  | (~\a[2]  ^ ~\a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[1]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  ^ \a[5] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[0]  | (\a[3]  ^ \a[4] ) | (~\a[2]  ^ ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[1]  | (~\a[2]  ^ ~\a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[2]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  ^ \a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n989_ = (~\a[8]  | ((~\b[0]  | (~\a[5]  ^ ~\a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[1]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  ^ \a[8] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )))) ^ ((~\b[1]  | (~\a[5]  ^ ~\a[6] ) | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] )) & (~\b[2]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  ^ \a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (\a[6]  ^ \a[7] ) | (~\a[5]  ^ ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )));
  assign new_n990_ = \a[5]  ^ (new_n991_ & (~new_n981_ | ((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))))));
  assign new_n991_ = (~\b[9]  | (~\a[2]  ^ ~\a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[10]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[8]  | (\a[3]  ^ \a[4] ) | (~\a[2]  ^ ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ));
  assign new_n992_ = \a[5]  ^ ((~\b[7]  | (\a[2]  ^ \a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[8]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[6]  | (\a[3]  ^ \a[4] ) | (\a[2]  ^ \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & ((\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n79_ & (~\b[7]  ^ \b[8] ))));
  assign new_n993_ = ~new_n968_ ^ (new_n863_ ^ ~new_n967_);
  assign new_n994_ = ~new_n965_ ^ (new_n877_ ^ ((~new_n880_ & (new_n782_ | (~new_n781_ & new_n789_) | (new_n781_ & ~new_n789_)) & (~new_n782_ | (~new_n781_ ^ new_n789_))) | (~new_n863_ & (new_n880_ | (~new_n782_ & (new_n781_ | ~new_n789_) & (~new_n781_ | new_n789_)) | (new_n782_ & (new_n781_ ^ new_n789_))) & (~new_n880_ | (~new_n782_ ^ (~new_n781_ ^ new_n789_))))));
  assign new_n995_ = \a[5]  ^ ((~new_n133_ | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[12]  | (\a[2]  ^ \a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[13]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[11]  | (\a[3]  ^ \a[4] ) | (\a[2]  ^ \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n996_ = new_n960_ & (~new_n882_ ^ (new_n855_ | (~new_n858_ & new_n881_)));
  assign new_n997_ = \a[5]  ^ ((~new_n186_ | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[15]  | (\a[2]  ^ \a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[16]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[14]  | (\a[3]  ^ \a[4] ) | (\a[2]  ^ \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n998_ = \a[5]  ^ ((~\b[13]  | (\a[2]  ^ \a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[14]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[12]  | (\a[3]  ^ \a[4] ) | (\a[2]  ^ \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & ((\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n142_ & (~\b[13]  ^ \b[14] ))));
  assign new_n999_ = ~new_n956_ ^ (new_n850_ ^ ~new_n955_);
  assign new_n1000_ = ~new_n953_ ^ ((~new_n848_ & ~new_n884_) ^ ((~new_n886_ & (new_n771_ | ~new_n794_) & (~new_n771_ | new_n794_)) | (~new_n850_ & (new_n886_ | (~new_n771_ & new_n794_) | (new_n771_ & ~new_n794_)) & (~new_n886_ | (~new_n771_ ^ new_n794_)))));
  assign new_n1001_ = \a[5]  ^ ((~new_n253_ | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & (~\b[18]  | (\a[2]  ^ \a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[19]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  ^ \a[5] )) & (~\b[17]  | (\a[3]  ^ \a[4] ) | (\a[2]  ^ \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n1002_ = new_n948_ & (~new_n888_ ^ (new_n843_ | (~new_n846_ & new_n887_)));
  assign new_n1003_ = \a[5]  ^ (((\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~new_n201_ ^ ~\b[19] )) & (~\b[19]  | (\a[2]  ^ \a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[18]  | (\a[3]  ^ \a[4] ) | (\a[2]  ^ \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n1004_ = \a[8]  ^ ((~new_n745_ ^ \a[11] ) ^ ((new_n746_ & \a[11] ) | (~new_n747_ & (new_n746_ | \a[11] ) & (~new_n746_ | ~\a[11] ))));
  assign new_n1005_ = \a[5]  ^ ((new_n823_ ^ \a[8] ) ^ (new_n824_ | (~new_n826_ & new_n891_)));
  assign new_n1006_ = new_n1008_ ^ (~new_n1007_ ^ ((~\a[11]  | (~new_n65_ & new_n899_) | (new_n65_ & ~new_n899_)) & (((~new_n894_ | ~\a[11] ) & ((new_n894_ & \a[11] ) | (~new_n894_ & ~\a[11] ) | ((~new_n897_ | ~\a[11] ) & (new_n898_ | (new_n897_ & \a[11] ) | (~new_n897_ & ~\a[11] ))))) | (\a[11]  & (new_n65_ | ~new_n899_) & (~new_n65_ | new_n899_)) | (~\a[11]  & (new_n65_ ^ new_n899_)))));
  assign new_n1007_ = (~new_n544_ | ~\a[20] ) & ((~new_n544_ & ~\a[20] ) | (new_n544_ & \a[20] ) | ((~new_n560_ | ~\a[20] ) & (new_n67_ | (new_n560_ & \a[20] ) | (~new_n560_ & ~\a[20] ))));
  assign new_n1008_ = ~new_n1009_ ^ (\a[17]  ^ (\a[29]  ^ \a[32] ));
  assign new_n1009_ = (~\a[35]  | (new_n553_ & new_n555_) | (~new_n553_ & ~new_n555_)) & (((~new_n549_ | ~\a[35] ) & ((new_n549_ & \a[35] ) | (~new_n549_ & ~\a[35] ) | ((~new_n540_ | ~\a[35] ) & (new_n548_ | (new_n540_ & \a[35] ) | (~new_n540_ & ~\a[35] ))))) | (\a[35]  & (~new_n553_ | ~new_n555_) & (new_n553_ | new_n555_)) | (~\a[35]  & (~new_n553_ ^ new_n555_)));
  assign new_n1010_ = (~\a[2]  | (~new_n908_ & (new_n907_ | \a[5] ) & (~new_n907_ | ~\a[5] )) | (new_n908_ & (new_n907_ ^ ~\a[5] ))) & (((~new_n1011_ | ~\a[2] ) & ((~new_n1011_ & ~\a[2] ) | (new_n1011_ & \a[2] ) | ((~new_n1012_ | ~\a[2] ) & (new_n1013_ | (new_n1012_ & \a[2] ) | (~new_n1012_ & ~\a[2] ))))) | (\a[2]  & (new_n908_ | (~new_n907_ & ~\a[5] ) | (new_n907_ & \a[5] )) & (~new_n908_ | (~new_n907_ ^ ~\a[5] ))) | (~\a[2]  & (new_n908_ ^ (~new_n907_ ^ ~\a[5] ))));
  assign new_n1011_ = ((\a[5]  & (new_n640_ | ~new_n911_) & (~new_n640_ | new_n911_)) | (((new_n913_ & \a[5] ) | ((~new_n913_ | ~\a[5] ) & (new_n913_ | \a[5] ) & ((new_n914_ & \a[5] ) | (~new_n915_ & (~new_n914_ | ~\a[5] ) & (new_n914_ | \a[5] ))))) & (~\a[5]  | (~new_n640_ & new_n911_) | (new_n640_ & ~new_n911_)) & (\a[5]  | (~new_n640_ ^ new_n911_)))) ^ (\a[5]  ^ (new_n912_ ^ (new_n909_ | (~new_n640_ & new_n911_))));
  assign new_n1012_ = ((new_n913_ & \a[5] ) | ((new_n913_ | \a[5] ) & (~new_n913_ | ~\a[5] ) & ((new_n914_ & \a[5] ) | (~new_n915_ & (~new_n914_ | ~\a[5] ) & (new_n914_ | \a[5] ))))) ^ (\a[5]  ^ (new_n640_ ^ ~new_n911_));
  assign new_n1013_ = (~\a[2]  | ((~new_n913_ | ~\a[5] ) & (new_n913_ | \a[5] ) & ((new_n914_ & \a[5] ) | (~new_n915_ & (~new_n914_ | ~\a[5] ) & (new_n914_ | \a[5] )))) | ((~new_n913_ ^ \a[5] ) & (~new_n914_ | ~\a[5] ) & (new_n915_ | (new_n914_ & \a[5] ) | (~new_n914_ & ~\a[5] )))) & (((~\a[2]  | (~new_n915_ & (~new_n914_ | ~\a[5] ) & (new_n914_ | \a[5] )) | (new_n915_ & (~new_n914_ ^ \a[5] ))) & (((~new_n1014_ | ~\a[2] ) & (((~new_n1015_ | ~\a[2] ) & (new_n1016_ | (~new_n1015_ & ~\a[2] ) | (new_n1015_ & \a[2] ))) | (new_n1014_ & \a[2] ) | (~new_n1014_ & ~\a[2] ))) | (\a[2]  & (new_n915_ | (new_n914_ & \a[5] ) | (~new_n914_ & ~\a[5] )) & (~new_n915_ | (new_n914_ ^ \a[5] ))) | (~\a[2]  & (new_n915_ ^ (new_n914_ ^ \a[5] ))))) | (\a[2]  & ((new_n913_ & \a[5] ) | (~new_n913_ & ~\a[5] ) | ((~new_n914_ | ~\a[5] ) & (new_n915_ | (new_n914_ & \a[5] ) | (~new_n914_ & ~\a[5] )))) & ((new_n913_ ^ \a[5] ) | (new_n914_ & \a[5] ) | (~new_n915_ & (~new_n914_ | ~\a[5] ) & (new_n914_ | \a[5] )))) | (~\a[2]  & ((~new_n913_ ^ \a[5] ) ^ ((new_n914_ & \a[5] ) | (~new_n915_ & (~new_n914_ | ~\a[5] ) & (new_n914_ | \a[5] ))))));
  assign new_n1014_ = ((\a[5]  & (new_n807_ | ~new_n917_) & (~new_n807_ | new_n917_)) | (((new_n919_ & \a[5] ) | ((~new_n919_ | ~\a[5] ) & (new_n919_ | \a[5] ) & ((new_n920_ & \a[5] ) | (~new_n921_ & (~new_n920_ | ~\a[5] ) & (new_n920_ | \a[5] ))))) & (~\a[5]  | (~new_n807_ & new_n917_) | (new_n807_ & ~new_n917_)) & (\a[5]  | (~new_n807_ ^ new_n917_)))) ^ (\a[5]  ^ (new_n918_ ^ (new_n916_ | (~new_n807_ & new_n917_))));
  assign new_n1015_ = ((new_n919_ & \a[5] ) | ((new_n919_ | \a[5] ) & (~new_n919_ | ~\a[5] ) & ((new_n920_ & \a[5] ) | (~new_n921_ & (~new_n920_ | ~\a[5] ) & (new_n920_ | \a[5] ))))) ^ (\a[5]  ^ (new_n807_ ^ ~new_n917_));
  assign new_n1016_ = (~\a[2]  | ((~new_n919_ | ~\a[5] ) & (new_n919_ | \a[5] ) & ((new_n920_ & \a[5] ) | ((~new_n920_ | ~\a[5] ) & (new_n920_ | \a[5] ) & ((new_n1017_ & \a[5] ) | (~new_n1018_ & (~new_n1017_ | ~\a[5] ) & (new_n1017_ | \a[5] )))))) | ((~new_n919_ ^ \a[5] ) & (~new_n920_ | ~\a[5] ) & ((new_n920_ & \a[5] ) | (~new_n920_ & ~\a[5] ) | ((~new_n1017_ | ~\a[5] ) & (new_n1018_ | (new_n1017_ & \a[5] ) | (~new_n1017_ & ~\a[5] )))))) & (((~\a[2]  | ((~new_n920_ | ~\a[5] ) & (new_n920_ | \a[5] ) & ((new_n1017_ & \a[5] ) | (~new_n1018_ & (~new_n1017_ | ~\a[5] ) & (new_n1017_ | \a[5] )))) | ((~new_n920_ ^ \a[5] ) & (~new_n1017_ | ~\a[5] ) & (new_n1018_ | (new_n1017_ & \a[5] ) | (~new_n1017_ & ~\a[5] )))) & (((~\a[2]  | (~new_n1018_ & (~new_n1017_ | ~\a[5] ) & (new_n1017_ | \a[5] )) | (new_n1018_ & (~new_n1017_ ^ \a[5] ))) & (((~new_n1019_ | ~\a[2] ) & (new_n1020_ | (~new_n1019_ & ~\a[2] ) | (new_n1019_ & \a[2] ))) | (\a[2]  & (new_n1018_ | (new_n1017_ & \a[5] ) | (~new_n1017_ & ~\a[5] )) & (~new_n1018_ | (new_n1017_ ^ \a[5] ))) | (~\a[2]  & (new_n1018_ ^ (new_n1017_ ^ \a[5] ))))) | (\a[2]  & ((new_n920_ & \a[5] ) | (~new_n920_ & ~\a[5] ) | ((~new_n1017_ | ~\a[5] ) & (new_n1018_ | (new_n1017_ & \a[5] ) | (~new_n1017_ & ~\a[5] )))) & ((new_n920_ ^ \a[5] ) | (new_n1017_ & \a[5] ) | (~new_n1018_ & (~new_n1017_ | ~\a[5] ) & (new_n1017_ | \a[5] )))) | (~\a[2]  & ((~new_n920_ ^ \a[5] ) ^ ((new_n1017_ & \a[5] ) | (~new_n1018_ & (~new_n1017_ | ~\a[5] ) & (new_n1017_ | \a[5] ))))))) | (\a[2]  & ((new_n919_ & \a[5] ) | (~new_n919_ & ~\a[5] ) | ((~new_n920_ | ~\a[5] ) & ((new_n920_ & \a[5] ) | (~new_n920_ & ~\a[5] ) | ((~new_n1017_ | ~\a[5] ) & (new_n1018_ | (new_n1017_ & \a[5] ) | (~new_n1017_ & ~\a[5] )))))) & ((new_n919_ ^ \a[5] ) | (new_n920_ & \a[5] ) | ((~new_n920_ | ~\a[5] ) & (new_n920_ | \a[5] ) & ((new_n1017_ & \a[5] ) | (~new_n1018_ & (~new_n1017_ | ~\a[5] ) & (new_n1017_ | \a[5] )))))) | (~\a[2]  & ((~new_n919_ ^ \a[5] ) ^ ((new_n920_ & \a[5] ) | ((~new_n920_ | ~\a[5] ) & (new_n920_ | \a[5] ) & ((new_n1017_ & \a[5] ) | (~new_n1018_ & (~new_n1017_ | ~\a[5] ) & (new_n1017_ | \a[5] ))))))));
  assign new_n1017_ = new_n810_ ^ ~new_n922_;
  assign new_n1018_ = (~new_n923_ | ~\a[5] ) & ((new_n923_ & \a[5] ) | (~new_n923_ & ~\a[5] ) | ((~new_n924_ | ~\a[5] ) & ((~new_n924_ & ~\a[5] ) | (new_n924_ & \a[5] ) | ((~new_n925_ | ~\a[5] ) & (new_n926_ | (new_n925_ & \a[5] ) | (~new_n925_ & ~\a[5] ))))));
  assign new_n1019_ = (new_n923_ ^ \a[5] ) ^ ((new_n924_ & \a[5] ) | ((new_n924_ | \a[5] ) & (~new_n924_ | ~\a[5] ) & ((new_n925_ & \a[5] ) | (~new_n926_ & (~new_n925_ | ~\a[5] ) & (new_n925_ | \a[5] )))));
  assign new_n1020_ = (~\a[2]  | ((~new_n924_ | ~\a[5] ) & (new_n924_ | \a[5] ) & ((new_n925_ & \a[5] ) | (~new_n926_ & (~new_n925_ | ~\a[5] ) & (new_n925_ | \a[5] )))) | ((~new_n924_ ^ \a[5] ) & (~new_n925_ | ~\a[5] ) & (new_n926_ | (new_n925_ & \a[5] ) | (~new_n925_ & ~\a[5] )))) & (((~\a[2]  | (~new_n926_ & (~new_n925_ | ~\a[5] ) & (new_n925_ | \a[5] )) | (new_n926_ & (~new_n925_ ^ \a[5] ))) & (((~new_n1021_ | ~\a[2] ) & (((~new_n1022_ | ~\a[2] ) & (new_n1024_ | (~new_n1022_ & ~\a[2] ) | (new_n1022_ & \a[2] ))) | (new_n1021_ & \a[2] ) | (~new_n1021_ & ~\a[2] ))) | (\a[2]  & (new_n926_ | (new_n925_ & \a[5] ) | (~new_n925_ & ~\a[5] )) & (~new_n926_ | (new_n925_ ^ \a[5] ))) | (~\a[2]  & (new_n926_ ^ (new_n925_ ^ \a[5] ))))) | (\a[2]  & ((new_n924_ & \a[5] ) | (~new_n924_ & ~\a[5] ) | ((~new_n925_ | ~\a[5] ) & (new_n926_ | (new_n925_ & \a[5] ) | (~new_n925_ & ~\a[5] )))) & ((new_n924_ ^ \a[5] ) | (new_n925_ & \a[5] ) | (~new_n926_ & (~new_n925_ | ~\a[5] ) & (new_n925_ | \a[5] )))) | (~\a[2]  & ((~new_n924_ ^ \a[5] ) ^ ((new_n925_ & \a[5] ) | (~new_n926_ & (~new_n925_ | ~\a[5] ) & (new_n925_ | \a[5] ))))));
  assign new_n1021_ = ((new_n927_ & \a[5] ) | ((~new_n927_ | ~\a[5] ) & (new_n927_ | \a[5] ) & ((new_n928_ & \a[5] ) | (((new_n929_ & \a[5] ) | (~new_n930_ & (new_n929_ | \a[5] ) & (~new_n929_ | ~\a[5] ))) & (~new_n928_ | ~\a[5] ) & (new_n928_ | \a[5] ))))) ^ (\a[5]  ^ (~new_n817_ ^ (new_n816_ ^ \a[8] )));
  assign new_n1022_ = (new_n927_ ^ \a[5] ) ^ ((new_n928_ & \a[5] ) | ((~new_n928_ | ~\a[5] ) & (new_n928_ | \a[5] ) & ((~new_n930_ & new_n1023_) | (new_n929_ & \a[5] ))));
  assign new_n1023_ = \a[5]  ^ ((new_n819_ ^ \a[8] ) ^ (new_n820_ | (~new_n821_ & new_n892_)));
  assign new_n1024_ = (~\a[2]  | ((~new_n928_ | ~\a[5] ) & (new_n928_ | \a[5] ) & ((new_n929_ & \a[5] ) | (~new_n930_ & (~new_n929_ | ~\a[5] ) & (new_n929_ | \a[5] )))) | ((~new_n928_ ^ \a[5] ) & (~new_n929_ | ~\a[5] ) & (new_n930_ | (new_n929_ & \a[5] ) | (~new_n929_ & ~\a[5] )))) & (((~\a[2]  | (~new_n930_ & (~new_n929_ | ~\a[5] ) & (new_n929_ | \a[5] )) | (new_n930_ & (~new_n929_ ^ \a[5] ))) & (((~new_n1025_ | ~\a[2] ) & (((~new_n1026_ | ~\a[2] ) & (new_n1028_ | (~new_n1026_ & ~\a[2] ) | (new_n1026_ & \a[2] ))) | (new_n1025_ & \a[2] ) | (~new_n1025_ & ~\a[2] ))) | (\a[2]  & (new_n930_ | (new_n929_ & \a[5] ) | (~new_n929_ & ~\a[5] )) & (~new_n930_ | (new_n929_ ^ \a[5] ))) | (~\a[2]  & (new_n930_ ^ (new_n929_ ^ \a[5] ))))) | (\a[2]  & ((new_n928_ & \a[5] ) | (~new_n928_ & ~\a[5] ) | ((~new_n929_ | ~\a[5] ) & (new_n930_ | (new_n929_ & \a[5] ) | (~new_n929_ & ~\a[5] )))) & ((new_n928_ ^ \a[5] ) | (new_n929_ & \a[5] ) | (~new_n930_ & (~new_n929_ | ~\a[5] ) & (new_n929_ | \a[5] )))) | (~\a[2]  & ((~new_n928_ ^ \a[5] ) ^ ((new_n929_ & \a[5] ) | (~new_n930_ & (~new_n929_ | ~\a[5] ) & (new_n929_ | \a[5] ))))));
  assign new_n1025_ = (\a[5]  ^ (new_n821_ ^ ~new_n892_)) ^ ((new_n931_ & \a[5] ) | ((~new_n931_ | ~\a[5] ) & (new_n931_ | \a[5] ) & ((new_n932_ & \a[5] ) | ((~new_n932_ | ~\a[5] ) & (new_n932_ | \a[5] ) & (new_n933_ | (~new_n934_ & new_n1005_))))));
  assign new_n1026_ = (~new_n931_ ^ ~\a[5] ) ^ ((new_n932_ & \a[5] ) | (new_n1027_ & (new_n933_ | (~new_n934_ & new_n1005_))));
  assign new_n1027_ = \a[5]  ^ ((~new_n822_ ^ ~\a[8] ) ^ ((new_n823_ & \a[8] ) | ((~new_n823_ | ~\a[8] ) & (new_n823_ | \a[8] ) & (new_n824_ | (~new_n826_ & new_n891_)))));
  assign new_n1028_ = (~\a[2]  | (new_n1027_ & (new_n933_ | (~new_n934_ & new_n1005_))) | (~new_n1027_ & ~new_n933_ & (new_n934_ | ~new_n1005_))) & (((~\a[2]  | (~new_n934_ & new_n1005_) | (new_n934_ & ~new_n1005_)) & (((~new_n1029_ | ~\a[2] ) & ((new_n1029_ & \a[2] ) | (~new_n1029_ & ~\a[2] ) | ((~new_n1030_ | ~\a[2] ) & (new_n1031_ | (new_n1030_ & \a[2] ) | (~new_n1030_ & ~\a[2] ))))) | (\a[2]  & (new_n934_ | ~new_n1005_) & (~new_n934_ | new_n1005_)) | (~\a[2]  & (new_n934_ ^ new_n1005_)))) | (\a[2]  & (~new_n1027_ | (~new_n933_ & (new_n934_ | ~new_n1005_))) & (new_n1027_ | new_n933_ | (~new_n934_ & new_n1005_))) | (~\a[2]  & (~new_n1027_ ^ (new_n933_ | (~new_n934_ & new_n1005_)))));
  assign new_n1029_ = (\a[5]  ^ (new_n826_ ^ ~new_n891_)) ^ ((new_n935_ & \a[5] ) | ((~new_n935_ | ~\a[5] ) & (new_n935_ | \a[5] ) & ((new_n936_ & \a[5] ) | ((~new_n936_ | ~\a[5] ) & (new_n936_ | \a[5] ) & ((\a[5]  & (new_n829_ | ~new_n1004_) & (~new_n829_ | new_n1004_)) | (~new_n937_ & (~\a[5]  | (~new_n829_ & new_n1004_) | (new_n829_ & ~new_n1004_)) & (\a[5]  | (~new_n829_ ^ new_n1004_))))))));
  assign new_n1030_ = ((new_n936_ & \a[5] ) | ((~new_n936_ | ~\a[5] ) & (new_n936_ | \a[5] ) & ((\a[5]  & (new_n829_ | ~new_n1004_) & (~new_n829_ | new_n1004_)) | (~new_n937_ & (~\a[5]  | (~new_n829_ & new_n1004_) | (new_n829_ & ~new_n1004_)) & (\a[5]  | (~new_n829_ ^ new_n1004_)))))) ^ (new_n935_ ^ \a[5] );
  assign new_n1031_ = (~\a[2]  | ((new_n1035_ | (new_n1096_ ^ ~\a[2] )) & ~new_n1096_ & ~new_n1097_ & (new_n937_ ^ new_n1033_))) & ((new_n1034_ & (new_n1032_ | (~new_n937_ & new_n1033_))) | (~new_n1034_ & ~new_n1032_ & (new_n937_ | ~new_n1033_)) | (~\a[2]  & (~new_n1097_ | (~new_n937_ & new_n1033_) | (new_n937_ & ~new_n1033_) | new_n1035_ | (new_n1096_ ^ ~\a[2] ))));
  assign new_n1032_ = \a[5]  & (~new_n829_ | new_n1004_) & (new_n829_ | ~new_n1004_);
  assign new_n1033_ = \a[5]  ^ (new_n829_ ^ ~new_n1004_);
  assign new_n1034_ = \a[5]  ^ (((\a[8]  & (((~new_n746_ | ~\a[11] ) & (new_n747_ | (new_n746_ & \a[11] ) | (~new_n746_ & ~\a[11] ))) | (~new_n745_ & \a[11] ) | (new_n745_ & ~\a[11] )) & ((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] )) | (~new_n745_ ^ \a[11] ))) | (~new_n829_ & (~\a[8]  | (((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] ))) & (new_n745_ | ~\a[11] ) & (~new_n745_ | \a[11] )) | ((~new_n746_ | ~\a[11] ) & (new_n747_ | (new_n746_ & \a[11] ) | (~new_n746_ & ~\a[11] )) & (new_n745_ ^ \a[11] ))) & (\a[8]  | (((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] ))) ^ (~new_n745_ ^ \a[11] ))))) ^ (\a[8]  ^ ((new_n827_ ^ \a[11] ) ^ ((~new_n745_ & \a[11] ) | (((new_n746_ & \a[11] ) | (~new_n747_ & (~new_n746_ | ~\a[11] ) & (new_n746_ | \a[11] ))) & (new_n745_ | ~\a[11] ) & (~new_n745_ | \a[11] ))))));
  assign new_n1035_ = (~\a[2]  | (new_n940_ & ~new_n1036_) | (~new_n940_ & new_n1036_)) & (((~new_n1037_ | ~\a[2] ) & ((~new_n1037_ & ~\a[2] ) | (new_n1037_ & \a[2] ) | ((~new_n1038_ | ~\a[2] ) & (new_n1041_ | (new_n1038_ & \a[2] ) | (~new_n1038_ & ~\a[2] ))))) | (\a[2]  & (~new_n940_ | new_n1036_) & (new_n940_ | ~new_n1036_)) | (~\a[2]  & (~new_n940_ ^ ~new_n1036_)));
  assign new_n1036_ = \a[5]  ^ ((new_n831_ ^ \a[8] ) ^ ((new_n832_ & \a[8] ) | (~new_n833_ & (new_n832_ | \a[8] ) & (~new_n832_ | ~\a[8] ))));
  assign new_n1037_ = ((\a[5]  & (new_n941_ | (new_n834_ & \a[8] ) | (~new_n834_ & ~\a[8] )) & (~new_n941_ | (new_n834_ ^ \a[8] ))) | (((new_n942_ & \a[5] ) | ((~new_n942_ | ~\a[5] ) & (new_n942_ | \a[5] ) & ((new_n943_ & \a[5] ) | (~new_n945_ & (~new_n943_ | ~\a[5] ) & (new_n943_ | \a[5] ))))) & (~\a[5]  | (~new_n941_ & (~new_n834_ | ~\a[8] ) & (new_n834_ | \a[8] )) | (new_n941_ & (~new_n834_ ^ \a[8] ))) & (\a[5]  | (~new_n941_ ^ (new_n834_ ^ \a[8] ))))) ^ (\a[5]  ^ ((new_n832_ ^ \a[8] ) ^ ((new_n834_ & \a[8] ) | (~new_n941_ & (~new_n834_ | ~\a[8] ) & (new_n834_ | \a[8] )))));
  assign new_n1038_ = (new_n1039_ ^ \a[5] ) ^ ((new_n942_ & \a[5] ) | ((new_n942_ | \a[5] ) & (~new_n942_ | ~\a[5] ) & ((new_n943_ & \a[5] ) | (~new_n945_ & (~new_n943_ | ~\a[5] ) & (new_n943_ | \a[5] )))));
  assign new_n1039_ = new_n1040_ ^ (new_n835_ | (~new_n835_ & ~new_n837_ & ((~new_n890_ & (new_n759_ | ~new_n800_) & (~new_n759_ | new_n800_)) | (~new_n838_ & (new_n890_ | (~new_n759_ & new_n800_) | (new_n759_ & ~new_n800_)) & (~new_n890_ | (~new_n759_ ^ new_n800_))))));
  assign new_n1040_ = \a[8]  ^ ((new_n752_ ^ ~new_n802_) ^ (new_n754_ | (new_n801_ & (new_n756_ | (~new_n759_ & new_n800_)))));
  assign new_n1041_ = (~\a[2]  | ((~new_n942_ | ~\a[5] ) & (new_n942_ | \a[5] ) & ((new_n943_ & \a[5] ) | ((~new_n943_ | ~\a[5] ) & (new_n943_ | \a[5] ) & ((new_n946_ & \a[5] ) | (~new_n1042_ & (~new_n946_ | ~\a[5] ) & (new_n946_ | \a[5] )))))) | ((~new_n942_ ^ \a[5] ) & (~new_n943_ | ~\a[5] ) & ((new_n943_ & \a[5] ) | (~new_n943_ & ~\a[5] ) | ((~new_n946_ | ~\a[5] ) & (new_n1042_ | (new_n946_ & \a[5] ) | (~new_n946_ & ~\a[5] )))))) & (((~\a[2]  | ((~new_n943_ | ~\a[5] ) & (new_n943_ | \a[5] ) & ((new_n946_ & \a[5] ) | (~new_n1042_ & (~new_n946_ | ~\a[5] ) & (new_n946_ | \a[5] )))) | ((~new_n943_ ^ \a[5] ) & (~new_n946_ | ~\a[5] ) & (new_n1042_ | (new_n946_ & \a[5] ) | (~new_n946_ & ~\a[5] )))) & (((~\a[2]  | (~new_n1042_ & (~new_n946_ | ~\a[5] ) & (new_n946_ | \a[5] )) | (new_n1042_ & (~new_n946_ ^ \a[5] ))) & (((~new_n1043_ | ~\a[2] ) & (new_n1044_ | (new_n1043_ & \a[2] ) | (~new_n1043_ & ~\a[2] ))) | (\a[2]  & (new_n1042_ | (new_n946_ & \a[5] ) | (~new_n946_ & ~\a[5] )) & (~new_n1042_ | (new_n946_ ^ \a[5] ))) | (~\a[2]  & (new_n1042_ ^ (new_n946_ ^ \a[5] ))))) | (\a[2]  & ((new_n943_ & \a[5] ) | (~new_n943_ & ~\a[5] ) | ((~new_n946_ | ~\a[5] ) & (new_n1042_ | (new_n946_ & \a[5] ) | (~new_n946_ & ~\a[5] )))) & ((new_n943_ ^ \a[5] ) | (new_n946_ & \a[5] ) | (~new_n1042_ & (~new_n946_ | ~\a[5] ) & (new_n946_ | \a[5] )))) | (~\a[2]  & ((~new_n943_ ^ \a[5] ) ^ ((new_n946_ & \a[5] ) | (~new_n1042_ & (~new_n946_ | ~\a[5] ) & (new_n946_ | \a[5] ))))))) | (\a[2]  & ((new_n942_ & \a[5] ) | (~new_n942_ & ~\a[5] ) | ((~new_n943_ | ~\a[5] ) & ((new_n943_ & \a[5] ) | (~new_n943_ & ~\a[5] ) | ((~new_n946_ | ~\a[5] ) & (new_n1042_ | (new_n946_ & \a[5] ) | (~new_n946_ & ~\a[5] )))))) & ((new_n942_ ^ \a[5] ) | (new_n943_ & \a[5] ) | ((~new_n943_ | ~\a[5] ) & (new_n943_ | \a[5] ) & ((new_n946_ & \a[5] ) | (~new_n1042_ & (~new_n946_ | ~\a[5] ) & (new_n946_ | \a[5] )))))) | (~\a[2]  & ((~new_n942_ ^ \a[5] ) ^ ((new_n943_ & \a[5] ) | ((~new_n943_ | ~\a[5] ) & (new_n943_ | \a[5] ) & ((new_n946_ & \a[5] ) | (~new_n1042_ & (~new_n946_ | ~\a[5] ) & (new_n946_ | \a[5] ))))))));
  assign new_n1042_ = ~new_n947_ & (new_n947_ | new_n1002_ | ((new_n1003_ | (~new_n846_ & new_n887_) | (new_n846_ & ~new_n887_)) & (new_n949_ | (~new_n1003_ & (new_n846_ | ~new_n887_) & (~new_n846_ | new_n887_)) | (new_n1003_ & (new_n846_ ^ new_n887_)))));
  assign new_n1043_ = (~new_n947_ & ~new_n1002_) ^ ((~new_n1003_ & (new_n846_ | ~new_n887_) & (~new_n846_ | new_n887_)) | (~new_n949_ & (new_n1003_ | (~new_n846_ & new_n887_) | (new_n846_ & ~new_n887_)) & (~new_n1003_ | (~new_n846_ ^ new_n887_))));
  assign new_n1044_ = (~\a[2]  | (new_n949_ & ~new_n1045_) | (~new_n949_ & new_n1045_)) & ((\a[2]  & (~new_n949_ | new_n1045_) & (new_n949_ | ~new_n1045_)) | (~\a[2]  & (~new_n949_ ^ ~new_n1045_)) | ((~new_n1046_ | ~\a[2] ) & ((new_n1046_ & \a[2] ) | (~new_n1046_ & ~\a[2] ) | (~new_n1047_ & (new_n1049_ | ~new_n1095_)))));
  assign new_n1045_ = ~new_n1003_ ^ (new_n846_ ^ ~new_n887_);
  assign new_n1046_ = (new_n950_ ^ ~new_n1001_) ^ (new_n952_ | (new_n1000_ & (new_n954_ | (~new_n957_ & new_n999_))));
  assign new_n1047_ = ~new_n1048_ & (~new_n1000_ | (~new_n954_ & (new_n957_ | ~new_n999_))) & (new_n1000_ | new_n954_ | (~new_n957_ & new_n999_));
  assign new_n1048_ = \a[2]  ^ (~\b[19]  | ((new_n201_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (\a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ))));
  assign new_n1049_ = (new_n1093_ | (new_n957_ & ~new_n999_) | (~new_n957_ & new_n999_)) & (((~new_n1050_ | new_n1094_) & ((~new_n1052_ & (new_n1054_ | ~new_n1092_)) | (~new_n1050_ & new_n1094_) | (new_n1050_ & ~new_n1094_))) | (~new_n1093_ & (~new_n957_ | new_n999_) & (new_n957_ | ~new_n999_)) | (new_n1093_ & (~new_n957_ ^ ~new_n999_)));
  assign new_n1050_ = new_n1051_ ^ (new_n959_ | (((~new_n998_ & (new_n858_ | ~new_n881_) & (~new_n858_ | new_n881_)) | (~new_n961_ & (new_n998_ | (~new_n858_ & new_n881_) | (new_n858_ & ~new_n881_)) & (~new_n998_ | (~new_n858_ ^ new_n881_)))) & ~new_n959_ & ~new_n996_));
  assign new_n1051_ = ~new_n997_ ^ ((new_n853_ | (new_n882_ & (new_n855_ | (~new_n858_ & new_n881_)))) ^ (new_n851_ ^ ~new_n883_));
  assign new_n1052_ = ~new_n1053_ & (new_n959_ | new_n996_ | ((new_n998_ | (~new_n858_ & new_n881_) | (new_n858_ & ~new_n881_)) & (new_n961_ | (~new_n998_ & (new_n858_ | ~new_n881_) & (~new_n858_ | new_n881_)) | (new_n998_ & (new_n858_ ^ new_n881_))))) & ((~new_n959_ & ~new_n996_) | (~new_n998_ & (new_n858_ | ~new_n881_) & (~new_n858_ | new_n881_)) | (~new_n961_ & (new_n998_ | (~new_n858_ & new_n881_) | (new_n858_ & ~new_n881_)) & (~new_n998_ | (~new_n858_ ^ new_n881_))));
  assign new_n1053_ = \a[2]  ^ ((~new_n199_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[16]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[18]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[17]  | \a[0]  | ~\a[1] ));
  assign new_n1054_ = (new_n1090_ | (new_n961_ & ~new_n1055_) | (~new_n961_ & new_n1055_)) & (((~new_n1056_ | new_n1091_) & ((~new_n1057_ & (new_n1059_ | ~new_n1089_)) | (~new_n1056_ & new_n1091_) | (new_n1056_ & ~new_n1091_))) | (~new_n1090_ & (~new_n961_ | new_n1055_) & (new_n961_ | ~new_n1055_)) | (new_n1090_ & (~new_n961_ ^ ~new_n1055_)));
  assign new_n1055_ = ~new_n998_ ^ (new_n858_ ^ ~new_n881_);
  assign new_n1056_ = (new_n962_ ^ ~new_n995_) ^ (new_n964_ | (new_n994_ & (new_n966_ | (~new_n969_ & new_n993_))));
  assign new_n1057_ = ~new_n1058_ & (~new_n994_ | (~new_n966_ & (new_n969_ | ~new_n993_))) & (new_n994_ | new_n966_ | (~new_n969_ & new_n993_));
  assign new_n1058_ = \a[2]  ^ ((~\b[13]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[15]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[14]  | \a[0]  | ~\a[1] ) & (~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | ((~\b[14]  | ~\b[15] ) & (\b[14]  | \b[15] ) & ((\b[13]  & \b[14] ) | (~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )))) | ((~\b[14]  ^ \b[15] ) & (~\b[13]  | ~\b[14] ) & (new_n142_ | (\b[13]  & \b[14] ) | (~\b[13]  & ~\b[14] )))));
  assign new_n1059_ = (new_n1087_ | (new_n969_ & ~new_n993_) | (~new_n969_ & new_n993_)) & (((~new_n1060_ | new_n1088_) & ((~new_n1062_ & (new_n1064_ | ~new_n1086_)) | (~new_n1060_ & new_n1088_) | (new_n1060_ & ~new_n1088_))) | (~new_n1087_ & (~new_n969_ | new_n993_) & (new_n969_ | ~new_n993_)) | (new_n1087_ & (~new_n969_ ^ ~new_n993_)));
  assign new_n1060_ = new_n1061_ ^ (new_n972_ | (new_n974_ & ((~new_n992_ & (new_n869_ | (~new_n868_ & new_n876_) | (new_n868_ & ~new_n876_)) & (~new_n869_ | (~new_n868_ ^ new_n876_))) | (~new_n975_ & (new_n992_ | (~new_n869_ & (new_n868_ | ~new_n876_) & (~new_n868_ | new_n876_)) | (new_n869_ & (new_n868_ ^ new_n876_))) & (~new_n992_ | (~new_n869_ ^ (~new_n868_ ^ new_n876_)))))));
  assign new_n1061_ = ~new_n990_ ^ ((new_n864_ ^ ~new_n865_) ^ ((new_n866_ & ~new_n867_) | ((~new_n866_ | new_n867_) & (new_n866_ | ~new_n867_) & ((~new_n868_ & new_n876_) | (~new_n869_ & (new_n868_ | ~new_n876_) & (~new_n868_ | new_n876_))))));
  assign new_n1062_ = ~new_n1063_ & (~new_n974_ | ((new_n992_ | (~new_n869_ & (new_n868_ | ~new_n876_) & (~new_n868_ | new_n876_)) | (new_n869_ & (new_n868_ ^ new_n876_))) & (new_n975_ | (~new_n992_ & (new_n869_ | (~new_n868_ & new_n876_) | (new_n868_ & ~new_n876_)) & (~new_n869_ | (~new_n868_ ^ new_n876_))) | (new_n992_ & (new_n869_ ^ (~new_n868_ ^ new_n876_)))))) & (new_n974_ | (~new_n992_ & (new_n869_ | (~new_n868_ & new_n876_) | (new_n868_ & ~new_n876_)) & (~new_n869_ | (~new_n868_ ^ new_n876_))) | (~new_n975_ & (new_n992_ | (~new_n869_ & (new_n868_ | ~new_n876_) & (~new_n868_ | new_n876_)) | (new_n869_ & (new_n868_ ^ new_n876_))) & (~new_n992_ | (~new_n869_ ^ (~new_n868_ ^ new_n876_)))));
  assign new_n1063_ = \a[2]  ^ ((~new_n107_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[10]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[12]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[11]  | \a[0]  | ~\a[1] ));
  assign new_n1064_ = (new_n1066_ | (new_n975_ & ~new_n1065_) | (~new_n975_ & new_n1065_)) & ((~new_n1066_ & (~new_n975_ | new_n1065_) & (new_n975_ | ~new_n1065_)) | (new_n1066_ & (~new_n975_ ^ ~new_n1065_)) | ((~new_n1067_ | new_n1085_) & ((~new_n1068_ & (new_n1070_ | ~new_n1084_)) | (~new_n1067_ & new_n1085_) | (new_n1067_ & ~new_n1085_))));
  assign new_n1065_ = ~new_n992_ ^ (~new_n869_ ^ (~new_n868_ ^ new_n876_));
  assign new_n1066_ = \a[2]  ^ ((~new_n135_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[9]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[11]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[10]  | \a[0]  | ~\a[1] ));
  assign new_n1067_ = (new_n976_ ^ ~new_n977_) ^ ((new_n978_ & ~new_n979_) | (((~new_n980_ & new_n989_) | (~new_n983_ & (new_n980_ | ~new_n989_) & (~new_n980_ | new_n989_))) & (~new_n978_ | new_n979_) & (new_n978_ | ~new_n979_)));
  assign new_n1068_ = ~new_n1069_ & ((new_n978_ & ~new_n979_) | (~new_n978_ & new_n979_) | ((new_n980_ | ~new_n989_) & (new_n983_ | (~new_n980_ & new_n989_) | (new_n980_ & ~new_n989_)))) & ((new_n978_ ^ ~new_n979_) | (~new_n980_ & new_n989_) | (~new_n983_ & (new_n980_ | ~new_n989_) & (~new_n980_ | new_n989_)));
  assign new_n1069_ = \a[2]  ^ ((~\b[7]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[9]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[8]  | \a[0]  | ~\a[1] ) & (~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))));
  assign new_n1070_ = (new_n1072_ | (new_n983_ & ~new_n1071_) | (~new_n983_ & new_n1071_)) & ((~new_n1072_ & (~new_n983_ | new_n1071_) & (new_n983_ | ~new_n1071_)) | (new_n1072_ & (~new_n983_ ^ ~new_n1071_)) | ((new_n1073_ | ~new_n1074_) & ((~new_n1073_ & new_n1074_) | (new_n1073_ & ~new_n1074_) | ((new_n1075_ | ~new_n1076_) & (new_n1077_ | (~new_n1075_ & new_n1076_) | (new_n1075_ & ~new_n1076_))))));
  assign new_n1071_ = new_n989_ ^ (~\a[5]  ^ (new_n982_ & (~new_n94_ | ~new_n981_)));
  assign new_n1072_ = \a[2]  ^ ((~\b[6]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[8]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[7]  | \a[0]  | ~\a[1] ) & ((~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n79_ & (~\b[7]  ^ \b[8] )) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )));
  assign new_n1073_ = \a[2]  ^ ((~new_n88_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[5]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[7]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[6]  | \a[0]  | ~\a[1] ));
  assign new_n1074_ = (new_n986_ | (~new_n987_ & new_n988_)) ^ (new_n985_ ^ (~\a[5]  ^ (new_n984_ & (~new_n98_ | ~new_n981_))));
  assign new_n1075_ = \a[2]  ^ ((~new_n91_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[4]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[6]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[5]  | \a[0]  | ~\a[1] ));
  assign new_n1076_ = new_n987_ ^ ~new_n988_;
  assign new_n1077_ = (~new_n1080_ | (\a[2]  ^ (new_n1079_ & (~new_n94_ | ~new_n1078_)))) & ((new_n1080_ & (~\a[2]  ^ (new_n1079_ & (~new_n94_ | ~new_n1078_)))) | (~new_n1080_ & (~\a[2]  | ~new_n1079_ | (new_n94_ & new_n1078_)) & (\a[2]  | (new_n1079_ & (~new_n94_ | ~new_n1078_)))) | ((new_n1081_ | ~new_n1082_) & (new_n1083_ | (~new_n1081_ & new_n1082_) | (new_n1081_ & ~new_n1082_))));
  assign new_n1078_ = \a[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] );
  assign new_n1079_ = (~\b[3]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[5]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[4]  | \a[0]  | ~\a[1] );
  assign new_n1080_ = (~\a[5]  | ((~\b[0]  | (~\a[2]  ^ ~\a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[1]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  ^ \a[5] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )))) ^ ((~\b[1]  | (~\a[2]  ^ ~\a[3] ) | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] )) & (~\b[2]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  ^ \a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (\a[3]  ^ \a[4] ) | (~\a[2]  ^ ~\a[3] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] )));
  assign new_n1081_ = \a[2]  ^ ((~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )))) | ((~\b[3]  ^ \b[4] ) & (~\b[2]  | ~\b[3] ) & ((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[4]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[3]  | \a[0]  | ~\a[1] ));
  assign new_n1082_ = ((\b[0]  & (\a[2]  ^ ~\a[3] ) & (~\a[3]  | ~\a[4] ) & (\a[3]  | \a[4] )) | (\b[1]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (~\a[4]  ^ \a[5] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (~\a[4]  | ~\a[5] ) & (\a[4]  | \a[5] ))) ^ (\a[5]  & \b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ));
  assign new_n1083_ = (~\b[0]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  ^ ((((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[3]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[1]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] )))) & ((\b[0]  & (~\a[2]  | ~\a[3] ) & (\a[2]  | \a[3] ) & (~\a[2]  ^ ((((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[3]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[1]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] )))) | ((~\b[0]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] )) & (~\a[2]  | (((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )) & ((\b[2]  ^ \b[3] ) | (\b[1]  & (\b[0]  | \b[2] ))) & \a[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] )) | (\b[3]  & \a[0]  & (~\a[1]  ^ \a[2] )) | (\b[1]  & ~\a[0]  & ~\a[1]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] )) | (\b[2]  & ~\a[0]  & \a[1] )) & (\a[2]  | ((((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[3]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[1]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] )))) | (\b[2]  & \a[0]  & (~\a[1]  ^ \a[2] )) | (\b[1]  & ~\a[0]  & \a[1] ) | (\b[0]  & ~\a[0]  & ~\a[1]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] )) | ((~\b[2]  ^ (\b[0]  | ~\b[1] )) & \a[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] )) | (\b[0]  & ~\a[0]  & \a[1] ) | (\b[1]  & \a[0]  & (~\a[1]  ^ \a[2] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & \a[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] )) | ~\a[2]  | (\a[0]  & \b[0] ));
  assign new_n1084_ = ~new_n1069_ ^ ((new_n978_ ^ ~new_n979_) ^ ((~new_n980_ & new_n989_) | (~new_n983_ & (new_n980_ | ~new_n989_) & (~new_n980_ | new_n989_))));
  assign new_n1085_ = \a[2]  ^ ((((~\b[9]  | ~\b[10] ) & (\b[9]  | \b[10] ) & ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n79_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))))) | ((~\b[9]  ^ \b[10] ) & (~\b[8]  | ~\b[9] ) & ((\b[8]  & \b[9] ) | (~\b[8]  & ~\b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n79_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))))) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[8]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[10]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[9]  | \a[0]  | ~\a[1] ));
  assign new_n1086_ = ~new_n1063_ ^ (new_n974_ ^ ((~new_n992_ & (new_n869_ | (~new_n868_ & new_n876_) | (new_n868_ & ~new_n876_)) & (~new_n869_ | (~new_n868_ ^ new_n876_))) | (~new_n975_ & (new_n992_ | (~new_n869_ & (new_n868_ | ~new_n876_) & (~new_n868_ | new_n876_)) | (new_n869_ & (new_n868_ ^ new_n876_))) & (~new_n992_ | (~new_n869_ ^ (~new_n868_ ^ new_n876_))))));
  assign new_n1087_ = \a[2]  ^ ((~\b[12]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[14]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[13]  | \a[0]  | ~\a[1] ) & ((~new_n142_ & (~\b[13]  | ~\b[14] ) & (\b[13]  | \b[14] )) | (new_n142_ & (~\b[13]  ^ \b[14] )) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )));
  assign new_n1088_ = \a[2]  ^ ((~new_n133_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[11]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[13]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[12]  | \a[0]  | ~\a[1] ));
  assign new_n1089_ = ~new_n1058_ ^ (new_n994_ ^ (new_n966_ | (~new_n969_ & new_n993_)));
  assign new_n1090_ = \a[2]  ^ ((~new_n144_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[15]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[17]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[16]  | \a[0]  | ~\a[1] ));
  assign new_n1091_ = \a[2]  ^ ((~new_n186_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[14]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[16]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[15]  | \a[0]  | ~\a[1] ));
  assign new_n1092_ = ~new_n1053_ ^ ((~new_n959_ & ~new_n996_) ^ ((~new_n998_ & (new_n858_ | ~new_n881_) & (~new_n858_ | new_n881_)) | (~new_n961_ & (new_n998_ | (~new_n858_ & new_n881_) | (new_n858_ & ~new_n881_)) & (~new_n998_ | (~new_n858_ ^ new_n881_)))));
  assign new_n1093_ = \a[2]  ^ (((new_n201_ ^ \b[19] ) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[18]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[19]  | \a[0]  | ~\a[1] ));
  assign new_n1094_ = \a[2]  ^ ((~new_n253_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[17]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[19]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[18]  | \a[0]  | ~\a[1] ));
  assign new_n1095_ = ~new_n1048_ ^ (new_n1000_ ^ (new_n954_ | (~new_n957_ & new_n999_)));
  assign new_n1096_ = (\a[5]  ^ ((~new_n938_ ^ ~\a[8] ) ^ ((new_n831_ & \a[8] ) | ((~new_n831_ | ~\a[8] ) & (new_n831_ | \a[8] ) & ((new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] ))))))) ^ ((\a[5]  & ((new_n831_ & \a[8] ) | (~new_n831_ & ~\a[8] ) | ((~new_n832_ | ~\a[8] ) & (new_n833_ | (new_n832_ & \a[8] ) | (~new_n832_ & ~\a[8] )))) & ((new_n831_ ^ \a[8] ) | (new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] )))) | (~new_n940_ & (~\a[5]  | ((~new_n831_ | ~\a[8] ) & (new_n831_ | \a[8] ) & ((new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] )))) | ((~new_n831_ ^ \a[8] ) & (~new_n832_ | ~\a[8] ) & (new_n833_ | (new_n832_ & \a[8] ) | (~new_n832_ & ~\a[8] )))) & (\a[5]  | ((new_n831_ ^ \a[8] ) ^ ((new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] )))))));
  assign new_n1097_ = (new_n939_ ^ \a[5] ) ^ ((\a[5]  & ((new_n938_ & \a[8] ) | (~new_n938_ & ~\a[8] ) | ((~new_n831_ | ~\a[8] ) & ((new_n831_ & \a[8] ) | (~new_n831_ & ~\a[8] ) | ((~new_n832_ | ~\a[8] ) & (new_n833_ | (new_n832_ & \a[8] ) | (~new_n832_ & ~\a[8] )))))) & ((new_n938_ ^ \a[8] ) | (new_n831_ & \a[8] ) | ((~new_n831_ | ~\a[8] ) & (new_n831_ | \a[8] ) & ((new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] )))))) | ((~\a[5]  | ((~new_n938_ | ~\a[8] ) & (new_n938_ | \a[8] ) & ((new_n831_ & \a[8] ) | ((~new_n831_ | ~\a[8] ) & (new_n831_ | \a[8] ) & ((new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] )))))) | ((~new_n938_ ^ \a[8] ) & (~new_n831_ | ~\a[8] ) & ((new_n831_ & \a[8] ) | (~new_n831_ & ~\a[8] ) | ((~new_n832_ | ~\a[8] ) & (new_n833_ | (new_n832_ & \a[8] ) | (~new_n832_ & ~\a[8] )))))) & (\a[5]  | ((new_n938_ ^ \a[8] ) ^ ((new_n831_ & \a[8] ) | ((~new_n831_ | ~\a[8] ) & (new_n831_ | \a[8] ) & ((new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] ))))))) & ((\a[5]  & ((new_n831_ & \a[8] ) | (~new_n831_ & ~\a[8] ) | ((~new_n832_ | ~\a[8] ) & (new_n833_ | (new_n832_ & \a[8] ) | (~new_n832_ & ~\a[8] )))) & ((new_n831_ ^ \a[8] ) | (new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] )))) | (~new_n940_ & (~\a[5]  | ((~new_n831_ | ~\a[8] ) & (new_n831_ | \a[8] ) & ((new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] )))) | ((~new_n831_ ^ \a[8] ) & (~new_n832_ | ~\a[8] ) & (new_n833_ | (new_n832_ & \a[8] ) | (~new_n832_ & ~\a[8] )))) & (\a[5]  | ((new_n831_ ^ \a[8] ) ^ ((new_n832_ & \a[8] ) | (~new_n833_ & (~new_n832_ | ~\a[8] ) & (new_n832_ | \a[8] )))))))));
  assign new_n1098_ = ((new_n1011_ & \a[2] ) | ((new_n1011_ | \a[2] ) & (~new_n1011_ | ~\a[2] ) & ((new_n1012_ & \a[2] ) | (~new_n1013_ & (~new_n1012_ | ~\a[2] ) & (new_n1012_ | \a[2] ))))) ^ (\a[2]  ^ (~new_n908_ ^ (~new_n907_ ^ ~\a[5] )));
  assign new_n1099_ = ((new_n1011_ ^ ~\a[2] ) ^ ((new_n1012_ & \a[2] ) | (((new_n1100_ & \a[2] ) | (~new_n1101_ & (~new_n1100_ | ~\a[2] ) & (new_n1100_ | \a[2] ))) & (~new_n1012_ | ~\a[2] ) & (new_n1012_ | \a[2] )))) & (((~new_n1100_ | ~\a[2] ) & (new_n1101_ | (new_n1100_ & \a[2] ) | (~new_n1100_ & ~\a[2] ))) ^ (new_n1012_ ^ \a[2] )) & (new_n1101_ ^ (new_n1100_ ^ \a[2] )) & ~new_n1102_ & new_n1103_;
  assign new_n1100_ = (~new_n913_ ^ ~\a[5] ) ^ ((new_n914_ & \a[5] ) | (~new_n915_ & (new_n914_ | \a[5] ) & (~new_n914_ | ~\a[5] )));
  assign new_n1101_ = (~\a[2]  | (~new_n915_ & (new_n914_ | \a[5] ) & (~new_n914_ | ~\a[5] )) | (new_n915_ & (new_n914_ ^ ~\a[5] ))) & (((~new_n1014_ | ~\a[2] ) & ((~new_n1014_ & ~\a[2] ) | (new_n1014_ & \a[2] ) | ((~new_n1015_ | ~\a[2] ) & (new_n1016_ | (new_n1015_ & \a[2] ) | (~new_n1015_ & ~\a[2] ))))) | (\a[2]  & (new_n915_ | (~new_n914_ & ~\a[5] ) | (new_n914_ & \a[5] )) & (~new_n915_ | (~new_n914_ ^ ~\a[5] ))) | (~\a[2]  & (new_n915_ ^ (~new_n914_ ^ ~\a[5] ))));
  assign new_n1102_ = ((new_n1014_ & \a[2] ) | ((new_n1014_ | \a[2] ) & (~new_n1014_ | ~\a[2] ) & ((new_n1015_ & \a[2] ) | (~new_n1016_ & (~new_n1015_ | ~\a[2] ) & (new_n1015_ | \a[2] ))))) ^ (\a[2]  ^ (~new_n915_ ^ (~new_n914_ ^ ~\a[5] )));
  assign new_n1103_ = ((new_n1014_ ^ ~\a[2] ) ^ ((new_n1015_ & \a[2] ) | (((new_n1104_ & \a[2] ) | (~new_n1105_ & (~new_n1104_ | ~\a[2] ) & (new_n1104_ | \a[2] ))) & (~new_n1015_ | ~\a[2] ) & (new_n1015_ | \a[2] )))) & (((~new_n1104_ | ~\a[2] ) & (new_n1105_ | (new_n1104_ & \a[2] ) | (~new_n1104_ & ~\a[2] ))) ^ (new_n1015_ ^ \a[2] )) & (new_n1105_ ^ (new_n1104_ ^ \a[2] )) & ~new_n1106_ & new_n1107_;
  assign new_n1104_ = (~new_n919_ ^ ~\a[5] ) ^ ((new_n920_ & \a[5] ) | (~new_n921_ & (new_n920_ | \a[5] ) & (~new_n920_ | ~\a[5] )));
  assign new_n1105_ = (~\a[2]  | ((new_n920_ | \a[5] ) & (~new_n920_ | ~\a[5] ) & ((new_n1017_ & \a[5] ) | (~new_n1018_ & (~new_n1017_ | ~\a[5] ) & (new_n1017_ | \a[5] )))) | ((new_n920_ ^ ~\a[5] ) & (~new_n1017_ | ~\a[5] ) & (new_n1018_ | (new_n1017_ & \a[5] ) | (~new_n1017_ & ~\a[5] )))) & (((~\a[2]  | (~new_n1018_ & (~new_n1017_ | ~\a[5] ) & (new_n1017_ | \a[5] )) | (new_n1018_ & (~new_n1017_ ^ \a[5] ))) & (((~new_n1019_ | ~\a[2] ) & (new_n1020_ | (new_n1019_ & \a[2] ) | (~new_n1019_ & ~\a[2] ))) | (\a[2]  & (new_n1018_ | (new_n1017_ & \a[5] ) | (~new_n1017_ & ~\a[5] )) & (~new_n1018_ | (new_n1017_ ^ \a[5] ))) | (~\a[2]  & (new_n1018_ ^ (new_n1017_ ^ \a[5] ))))) | (\a[2]  & ((~new_n920_ & ~\a[5] ) | (new_n920_ & \a[5] ) | ((~new_n1017_ | ~\a[5] ) & (new_n1018_ | (new_n1017_ & \a[5] ) | (~new_n1017_ & ~\a[5] )))) & ((~new_n920_ ^ ~\a[5] ) | (new_n1017_ & \a[5] ) | (~new_n1018_ & (~new_n1017_ | ~\a[5] ) & (new_n1017_ | \a[5] )))) | (~\a[2]  & ((new_n920_ ^ ~\a[5] ) ^ ((new_n1017_ & \a[5] ) | (~new_n1018_ & (~new_n1017_ | ~\a[5] ) & (new_n1017_ | \a[5] ))))));
  assign new_n1106_ = ((\a[2]  & (new_n1018_ | (new_n1017_ & \a[5] ) | (~new_n1017_ & ~\a[5] )) & (~new_n1018_ | (new_n1017_ ^ \a[5] ))) | (((new_n1019_ & \a[2] ) | (~new_n1020_ & (~new_n1019_ | ~\a[2] ) & (new_n1019_ | \a[2] ))) & (~\a[2]  | (~new_n1018_ & (~new_n1017_ | ~\a[5] ) & (new_n1017_ | \a[5] )) | (new_n1018_ & (~new_n1017_ ^ \a[5] ))) & (\a[2]  | (~new_n1018_ ^ (new_n1017_ ^ \a[5] ))))) ^ (\a[2]  ^ ((~new_n920_ ^ ~\a[5] ) ^ ((new_n1017_ & \a[5] ) | (~new_n1018_ & (~new_n1017_ | ~\a[5] ) & (new_n1017_ | \a[5] )))));
  assign new_n1107_ = ((~new_n1108_ ^ \a[2] ) ^ ((new_n1019_ & \a[2] ) | ((~new_n1019_ | ~\a[2] ) & (new_n1019_ | \a[2] ) & ((new_n1109_ & \a[2] ) | (~new_n1110_ & (new_n1109_ | \a[2] ) & (~new_n1109_ | ~\a[2] )))))) & ((~new_n1019_ ^ \a[2] ) ^ ((new_n1109_ & \a[2] ) | (~new_n1110_ & (new_n1109_ | \a[2] ) & (~new_n1109_ | ~\a[2] )))) & new_n1112_ & (new_n1110_ ^ (~new_n1109_ ^ ~\a[2] ));
  assign new_n1108_ = ((new_n923_ & \a[5] ) | ((~new_n923_ | ~\a[5] ) & (new_n923_ | \a[5] ) & ((new_n924_ & \a[5] ) | (((new_n925_ & \a[5] ) | (~new_n926_ & (new_n925_ | \a[5] ) & (~new_n925_ | ~\a[5] ))) & (~new_n924_ | ~\a[5] ) & (new_n924_ | \a[5] ))))) ^ (\a[5]  ^ (new_n810_ ^ ~new_n922_));
  assign new_n1109_ = (~new_n924_ ^ ~\a[5] ) ^ ((new_n925_ & \a[5] ) | (~new_n926_ & (new_n925_ | \a[5] ) & (~new_n925_ | ~\a[5] )));
  assign new_n1110_ = (~\a[2]  | (new_n926_ & ~new_n1111_) | (~new_n926_ & new_n1111_)) & (((~new_n1021_ | ~\a[2] ) & ((~new_n1021_ & ~\a[2] ) | (new_n1021_ & \a[2] ) | ((~new_n1022_ | ~\a[2] ) & (new_n1024_ | (new_n1022_ & \a[2] ) | (~new_n1022_ & ~\a[2] ))))) | (\a[2]  & (~new_n926_ | new_n1111_) & (new_n926_ | ~new_n1111_)) | (~\a[2]  & (~new_n926_ ^ ~new_n1111_)));
  assign new_n1111_ = \a[5]  ^ ((new_n815_ ^ \a[8] ) ^ ((new_n816_ & \a[8] ) | (~new_n817_ & (new_n816_ | \a[8] ) & (~new_n816_ | ~\a[8] ))));
  assign new_n1112_ = ((\a[2]  ^ (new_n926_ ^ ~new_n1111_)) ^ ((~new_n1021_ | ~\a[2] ) & ((new_n1021_ & \a[2] ) | (~new_n1021_ & ~\a[2] ) | ((~new_n1022_ | ~\a[2] ) & ((new_n1022_ & \a[2] ) | (~new_n1022_ & ~\a[2] ) | ((~new_n1113_ | ~\a[2] ) & (new_n1114_ | (new_n1113_ & \a[2] ) | (~new_n1113_ & ~\a[2] )))))))) & ((~new_n1021_ ^ \a[2] ) ^ ((new_n1022_ & \a[2] ) | ((~new_n1022_ | ~\a[2] ) & (new_n1022_ | \a[2] ) & ((new_n1113_ & \a[2] ) | (~new_n1114_ & (~new_n1113_ | ~\a[2] ) & (new_n1113_ | \a[2] )))))) & ((~new_n1022_ ^ \a[2] ) ^ ((new_n1113_ & \a[2] ) | (~new_n1114_ & (~new_n1113_ | ~\a[2] ) & (new_n1113_ | \a[2] )))) & new_n1115_ & (new_n1114_ ^ (new_n1113_ ^ \a[2] ));
  assign new_n1113_ = (~new_n928_ ^ ~\a[5] ) ^ ((new_n929_ & \a[5] ) | (~new_n930_ & (new_n929_ | \a[5] ) & (~new_n929_ | ~\a[5] )));
  assign new_n1114_ = (~\a[2]  | (new_n930_ & ~new_n1023_) | (~new_n930_ & new_n1023_)) & (((~new_n1025_ | ~\a[2] ) & ((~new_n1025_ & ~\a[2] ) | (new_n1025_ & \a[2] ) | ((~new_n1026_ | ~\a[2] ) & (new_n1028_ | (new_n1026_ & \a[2] ) | (~new_n1026_ & ~\a[2] ))))) | (\a[2]  & (~new_n930_ | new_n1023_) & (new_n930_ | ~new_n1023_)) | (~\a[2]  & (~new_n930_ ^ ~new_n1023_)));
  assign new_n1115_ = ((\a[2]  ^ (new_n930_ ^ ~new_n1023_)) ^ ((~new_n1025_ | ~\a[2] ) & ((new_n1025_ & \a[2] ) | (~new_n1025_ & ~\a[2] ) | ((~new_n1026_ | ~\a[2] ) & ((new_n1026_ & \a[2] ) | (~new_n1026_ & ~\a[2] ) | ((~new_n1116_ | ~\a[2] ) & (new_n1117_ | (new_n1116_ & \a[2] ) | (~new_n1116_ & ~\a[2] )))))))) & ((~new_n1025_ ^ \a[2] ) ^ ((new_n1026_ & \a[2] ) | ((~new_n1026_ | ~\a[2] ) & (new_n1026_ | \a[2] ) & ((new_n1116_ & \a[2] ) | (~new_n1117_ & (~new_n1116_ | ~\a[2] ) & (new_n1116_ | \a[2] )))))) & ((new_n1026_ ^ \a[2] ) | (new_n1116_ & \a[2] ) | (~new_n1117_ & (~new_n1116_ | ~\a[2] ) & (new_n1116_ | \a[2] ))) & ((new_n1026_ & \a[2] ) | (~new_n1026_ & ~\a[2] ) | ((~new_n1116_ | ~\a[2] ) & (new_n1117_ | (new_n1116_ & \a[2] ) | (~new_n1116_ & ~\a[2] )))) & (~new_n1117_ | (new_n1116_ ^ \a[2] )) & new_n1118_ & (new_n1117_ | (new_n1116_ & \a[2] ) | (~new_n1116_ & ~\a[2] ));
  assign new_n1116_ = new_n1027_ ^ (new_n933_ | (~new_n934_ & new_n1005_));
  assign new_n1117_ = (~\a[2]  | (new_n934_ & ~new_n1005_) | (~new_n934_ & new_n1005_)) & (((~new_n1029_ | ~\a[2] ) & ((~new_n1029_ & ~\a[2] ) | (new_n1029_ & \a[2] ) | ((~new_n1030_ | ~\a[2] ) & (new_n1031_ | (new_n1030_ & \a[2] ) | (~new_n1030_ & ~\a[2] ))))) | (\a[2]  & (~new_n934_ | new_n1005_) & (new_n934_ | ~new_n1005_)) | (~\a[2]  & (~new_n934_ ^ ~new_n1005_)));
  assign new_n1118_ = ((new_n1029_ & \a[2] ) | ((~new_n1029_ | ~\a[2] ) & (new_n1029_ | \a[2] ) & ((new_n1030_ & \a[2] ) | (~new_n1031_ & (~new_n1030_ | ~\a[2] ) & (new_n1030_ | \a[2] )))) | (\a[2]  ^ (new_n934_ ^ ~new_n1005_))) & (((~new_n1029_ | ~\a[2] ) & ((new_n1029_ & \a[2] ) | (~new_n1029_ & ~\a[2] ) | ((~new_n1030_ | ~\a[2] ) & (new_n1031_ | (new_n1030_ & \a[2] ) | (~new_n1030_ & ~\a[2] ))))) | (\a[2]  & (~new_n934_ | new_n1005_) & (new_n934_ | ~new_n1005_)) | (~\a[2]  & (~new_n934_ ^ ~new_n1005_))) & ((~new_n1029_ ^ \a[2] ) ^ ((new_n1030_ & \a[2] ) | (~new_n1031_ & (~new_n1030_ | ~\a[2] ) & (new_n1030_ | \a[2] )))) & (~new_n1031_ | (new_n1030_ ^ \a[2] )) & (new_n1031_ | (new_n1030_ & \a[2] ) | (~new_n1030_ & ~\a[2] )) & new_n1119_ & new_n1166_;
  assign new_n1119_ = new_n1122_ & (new_n1120_ | ~new_n1121_) & (~new_n1120_ | new_n1121_) & (~new_n937_ ^ ~new_n1033_) & (new_n1097_ ^ (new_n1096_ | ~\a[2] ));
  assign new_n1120_ = (~new_n1037_ | ~\a[2] ) & ((~new_n1037_ & ~\a[2] ) | (new_n1037_ & \a[2] ) | ((~new_n1038_ | ~\a[2] ) & (new_n1041_ | (~new_n1038_ & ~\a[2] ) | (new_n1038_ & \a[2] ))));
  assign new_n1121_ = \a[2]  ^ (new_n940_ ^ ~new_n1036_);
  assign new_n1122_ = ((new_n1037_ ^ ~\a[2] ) ^ ((new_n1038_ & \a[2] ) | (~new_n1041_ & (~new_n1038_ | ~\a[2] ) & (new_n1038_ | \a[2] )))) & (~new_n1041_ | (new_n1038_ ^ \a[2] )) & new_n1128_ & (~new_n1123_ ^ ~new_n1127_) & (new_n1041_ | (new_n1038_ & \a[2] ) | (~new_n1038_ & ~\a[2] ));
  assign new_n1123_ = (~\a[2]  | (new_n945_ & ~new_n1124_) | (~new_n945_ & new_n1124_)) & (((~new_n1125_ | ~\a[2] ) & ((~new_n1125_ & ~\a[2] ) | (new_n1125_ & \a[2] ) | ((~new_n1043_ | ~\a[2] ) & (new_n1044_ | (new_n1043_ & \a[2] ) | (~new_n1043_ & ~\a[2] ))))) | (\a[2]  & (~new_n945_ | new_n1124_) & (new_n945_ | ~new_n1124_)) | (~\a[2]  & (~new_n945_ ^ ~new_n1124_)));
  assign new_n1124_ = \a[5]  ^ (new_n838_ ^ ~new_n944_);
  assign new_n1125_ = new_n1126_ ^ (new_n947_ | (((~new_n1003_ & (new_n846_ | ~new_n887_) & (~new_n846_ | new_n887_)) | (~new_n949_ & (new_n1003_ | (~new_n846_ & new_n887_) | (new_n846_ & ~new_n887_)) & (~new_n1003_ | (~new_n846_ ^ new_n887_)))) & ~new_n947_ & ~new_n1002_));
  assign new_n1126_ = \a[5]  ^ ((new_n839_ ^ ~new_n889_) ^ (new_n841_ | (new_n888_ & (new_n843_ | (~new_n846_ & new_n887_)))));
  assign new_n1127_ = \a[2]  ^ ((new_n942_ ^ \a[5] ) ^ ((new_n943_ & \a[5] ) | (~new_n945_ & (new_n943_ | \a[5] ) & (~new_n943_ | ~\a[5] ))));
  assign new_n1128_ = ((\a[2]  ^ (new_n945_ ^ ~new_n1124_)) | (new_n1125_ & \a[2] ) | ((~new_n1125_ | ~\a[2] ) & (new_n1125_ | \a[2] ) & ((new_n1043_ & \a[2] ) | ((~new_n1043_ | ~\a[2] ) & (new_n1043_ | \a[2] ) & ((new_n1129_ & \a[2] ) | (~new_n1130_ & (~new_n1129_ | ~\a[2] ) & (new_n1129_ | \a[2] ))))))) & ((\a[2]  & (~new_n945_ | new_n1124_) & (new_n945_ | ~new_n1124_)) | (~\a[2]  & (~new_n945_ ^ ~new_n1124_)) | ((~new_n1125_ | ~\a[2] ) & ((new_n1125_ & \a[2] ) | (~new_n1125_ & ~\a[2] ) | ((~new_n1043_ | ~\a[2] ) & ((new_n1043_ & \a[2] ) | (~new_n1043_ & ~\a[2] ) | ((~new_n1129_ | ~\a[2] ) & (new_n1130_ | (new_n1129_ & \a[2] ) | (~new_n1129_ & ~\a[2] )))))))) & ((~new_n1125_ ^ \a[2] ) ^ ((new_n1043_ & \a[2] ) | ((~new_n1043_ | ~\a[2] ) & (new_n1043_ | \a[2] ) & ((new_n1129_ & \a[2] ) | (~new_n1130_ & (~new_n1129_ | ~\a[2] ) & (new_n1129_ | \a[2] )))))) & ((~new_n1043_ ^ \a[2] ) ^ ((new_n1129_ & \a[2] ) | (~new_n1130_ & (~new_n1129_ | ~\a[2] ) & (new_n1129_ | \a[2] )))) & (~new_n1130_ | (new_n1129_ ^ \a[2] )) & new_n1131_ & (new_n1130_ | (new_n1129_ & \a[2] ) | (~new_n1129_ & ~\a[2] ));
  assign new_n1129_ = new_n949_ ^ ~new_n1045_;
  assign new_n1130_ = (~new_n1046_ | ~\a[2] ) & ((~new_n1047_ & (new_n1049_ | ~new_n1095_)) | (new_n1046_ & \a[2] ) | (~new_n1046_ & ~\a[2] ));
  assign new_n1131_ = (~new_n1133_ ^ (new_n1047_ | (new_n1095_ & ((~new_n1093_ & (new_n957_ | ~new_n999_) & (~new_n957_ | new_n999_)) | (~new_n1132_ & (new_n1093_ | (~new_n957_ & new_n999_) | (new_n957_ & ~new_n999_)) & (~new_n1093_ | (~new_n957_ ^ new_n999_))))))) & (~new_n1095_ ^ ((~new_n1093_ & (new_n957_ | ~new_n999_) & (~new_n957_ | new_n999_)) | (~new_n1132_ & (new_n1093_ | (~new_n957_ & new_n999_) | (new_n957_ & ~new_n999_)) & (~new_n1093_ | (~new_n957_ ^ new_n999_))))) & (~new_n1132_ | (~new_n1093_ ^ (~new_n957_ ^ new_n999_))) & new_n1134_ & (new_n1132_ | (~new_n1093_ & (new_n957_ | ~new_n999_) & (~new_n957_ | new_n999_)) | (new_n1093_ & (new_n957_ ^ new_n999_)));
  assign new_n1132_ = (~new_n1050_ | new_n1094_) & ((~new_n1052_ & (new_n1054_ | ~new_n1092_)) | (~new_n1050_ & new_n1094_) | (new_n1050_ & ~new_n1094_));
  assign new_n1133_ = \a[2]  ^ ((new_n950_ ^ ~new_n1001_) ^ (new_n952_ | (new_n1000_ & (new_n954_ | (~new_n957_ & new_n999_)))));
  assign new_n1134_ = ((~new_n1050_ ^ ~new_n1094_) ^ (new_n1052_ | (~new_n1054_ & new_n1092_))) & (~new_n1054_ | new_n1092_) & (new_n1054_ | ~new_n1092_) & new_n1137_ & (~new_n1135_ ^ ~new_n1136_);
  assign new_n1135_ = (~new_n1056_ | new_n1091_) & ((~new_n1057_ & (new_n1059_ | ~new_n1089_)) | (~new_n1056_ & new_n1091_) | (new_n1056_ & ~new_n1091_));
  assign new_n1136_ = ~new_n1090_ ^ (new_n961_ ^ ~new_n1055_);
  assign new_n1137_ = (new_n1141_ | new_n1057_ | (new_n1089_ & (new_n1138_ | (~new_n1139_ & ~new_n1138_ & ~new_n1140_)))) & (~new_n1141_ | (~new_n1057_ & (~new_n1089_ | (~new_n1138_ & (new_n1139_ | new_n1138_ | new_n1140_))))) & (new_n1089_ | new_n1138_ | (~new_n1139_ & ~new_n1138_ & ~new_n1140_)) & (~new_n1089_ | (~new_n1138_ & (new_n1139_ | new_n1138_ | new_n1140_))) & (~new_n1139_ | (~new_n1138_ & ~new_n1140_)) & ~new_n1142_ & new_n1143_ & (new_n1139_ | new_n1138_ | new_n1140_);
  assign new_n1138_ = ~new_n1087_ & (~new_n969_ | new_n993_) & (new_n969_ | ~new_n993_);
  assign new_n1139_ = (~new_n1060_ | new_n1088_) & ((~new_n1062_ & (new_n1064_ | ~new_n1086_)) | (~new_n1060_ & new_n1088_) | (new_n1060_ & ~new_n1088_));
  assign new_n1140_ = new_n1087_ & (~new_n969_ ^ ~new_n993_);
  assign new_n1141_ = ~new_n1091_ ^ ((new_n964_ | (new_n994_ & (new_n966_ | (~new_n969_ & new_n993_)))) ^ (new_n962_ ^ ~new_n995_));
  assign new_n1142_ = (new_n1062_ | (~new_n1064_ & new_n1086_)) ^ (~new_n1060_ ^ new_n1088_);
  assign new_n1143_ = (~new_n1086_ ^ (new_n1144_ | (~new_n1144_ & ~new_n1147_ & (new_n1145_ | (new_n1067_ & ~new_n1085_))))) & ((~new_n1144_ & ~new_n1147_) | new_n1145_ | (new_n1067_ & ~new_n1085_)) & (new_n1144_ | new_n1147_ | (~new_n1145_ & (~new_n1067_ | new_n1085_))) & ~new_n1148_ & ~new_n1145_ & new_n1149_;
  assign new_n1144_ = ~new_n1066_ & (~new_n975_ | new_n1065_) & (new_n975_ | ~new_n1065_);
  assign new_n1145_ = new_n1146_ & (new_n1068_ | (~new_n1070_ & new_n1084_));
  assign new_n1146_ = ~new_n1085_ ^ ((new_n976_ ^ ~new_n977_) ^ ((new_n978_ & ~new_n979_) | ((~new_n978_ | new_n979_) & (new_n978_ | ~new_n979_) & ((~new_n980_ & new_n989_) | (~new_n983_ & (new_n980_ | ~new_n989_) & (~new_n980_ | new_n989_))))));
  assign new_n1147_ = new_n1066_ & (~new_n975_ ^ ~new_n1065_);
  assign new_n1148_ = ~new_n1146_ & ~new_n1068_ & (new_n1070_ | ~new_n1084_);
  assign new_n1149_ = (~new_n1070_ ^ ~new_n1084_) & (new_n1151_ | new_n1150_ | (~new_n1073_ & new_n1074_)) & (~new_n1151_ | (~new_n1150_ & (new_n1073_ | ~new_n1074_))) & ~new_n1152_ & ~new_n1150_ & new_n1153_;
  assign new_n1150_ = (~new_n1073_ | new_n1074_) & (new_n1073_ | ~new_n1074_) & ((~new_n1075_ & new_n1076_) | (~new_n1077_ & (~new_n1075_ | new_n1076_) & (new_n1075_ | ~new_n1076_)));
  assign new_n1151_ = ~new_n1072_ ^ (new_n983_ ^ ~new_n1071_);
  assign new_n1152_ = (~new_n1073_ ^ ~new_n1074_) & (new_n1075_ | ~new_n1076_) & (new_n1077_ | (new_n1075_ & ~new_n1076_) | (~new_n1075_ & new_n1076_));
  assign new_n1153_ = (~new_n1077_ | (new_n1075_ ^ ~new_n1076_)) & (new_n1077_ | (new_n1075_ & ~new_n1076_) | (~new_n1075_ & new_n1076_)) & ~new_n1154_ & ~new_n1155_ & ~new_n1165_ & ~new_n1156_ & new_n1162_;
  assign new_n1154_ = (new_n1080_ ^ (~\a[2]  ^ (new_n1079_ & (~new_n94_ | ~new_n1078_)))) ^ ((~new_n1081_ & new_n1082_) | (~new_n1083_ & (new_n1081_ | ~new_n1082_) & (~new_n1081_ | new_n1082_)));
  assign new_n1155_ = ~new_n1083_ ^ (new_n1081_ ^ ~new_n1082_);
  assign new_n1156_ = new_n1157_ & new_n1158_ & new_n1159_ & new_n1160_ & new_n1161_;
  assign new_n1157_ = ~\a[27]  & ~\a[28]  & ~\a[25]  & ~\a[26]  & ~\a[15]  & ~\a[16]  & ~\a[30]  & ~\a[31] ;
  assign new_n1158_ = ~\a[17]  & ~\a[18]  & ~\a[19]  & ~\a[20]  & ~\a[21]  & ~\a[22]  & ~\a[23]  & ~\a[24] ;
  assign new_n1159_ = ~\a[29]  & ~\a[32]  & ~\a[37]  & ~\a[38]  & ~\a[35]  & ~\a[36] ;
  assign new_n1160_ = ~\a[1]  & ~\a[2]  & ~\a[3]  & ~\a[4]  & ~\a[7]  & ~\a[8]  & ~\a[33]  & ~\a[34] ;
  assign new_n1161_ = ~\a[5]  & ~\a[6]  & ~\a[9]  & ~\a[10]  & ~\a[11]  & ~\a[12]  & ~\a[13]  & ~\a[14] ;
  assign new_n1162_ = \a[0]  & \b[0]  & (~new_n1163_ | ~new_n1164_ | \b[19]  | \b[1]  | \b[2] );
  assign new_n1163_ = ~\b[11]  & ~\b[12]  & ~\b[13]  & ~\b[14]  & ~\b[15]  & ~\b[16]  & ~\b[17]  & ~\b[18] ;
  assign new_n1164_ = ~\b[3]  & ~\b[4]  & ~\b[5]  & ~\b[6]  & ~\b[7]  & ~\b[8]  & ~\b[9]  & ~\b[10] ;
  assign new_n1165_ = ((\b[0]  & (~\a[2]  | ~\a[3] ) & (\a[2]  | \a[3] )) ^ (~\a[2]  ^ ((((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[3]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[1]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] )))) ? ((\b[2]  & \a[0]  & (~\a[1]  ^ \a[2] )) | (\b[1]  & ~\a[0]  & \a[1] ) | (\b[0]  & ~\a[0]  & ~\a[1]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] )) | ((~\b[2]  ^ (\b[0]  | ~\b[1] )) & \a[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] )) | (\b[0]  & ~\a[0]  & \a[1] ) | (\b[1]  & \a[0]  & (~\a[1]  ^ \a[2] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & \a[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] )) | ~\a[2]  | (\a[0]  & \b[0] )) : ((\a[2]  & (~\a[0]  | ~\b[0]  | ((~\b[1]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ))))) | (((~\b[2]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[1]  | \a[0]  | ~\a[1] ) & (~\b[0]  | \a[0]  | \a[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & ((\b[2]  ^ (\b[0]  | ~\b[1] )) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ))) ? ((\b[0]  & ~\a[0]  & \a[1] ) | (\b[1]  & \a[0]  & (~\a[1]  ^ \a[2] )) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & \a[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] ))) : ~\a[2] ));
  assign new_n1166_ = (~new_n1035_ | (~new_n1096_ & \a[2] ) | (new_n1096_ & ~\a[2] )) & (~new_n1034_ ^ (new_n1032_ | (~new_n937_ & new_n1033_))) & (new_n1035_ | (~new_n1096_ ^ \a[2] ));
  assign new_n1167_ = (~\a[11]  ^ \a[14] ) ^ ((~\a[17]  | ((~new_n544_ ^ \a[20] ) & (~new_n560_ | ~\a[20] ) & (new_n67_ | (new_n560_ & \a[20] ) | (~new_n560_ & ~\a[20] ))) | ((~new_n544_ | ~\a[20] ) & (new_n544_ | \a[20] ) & ((new_n560_ & \a[20] ) | (~new_n67_ & (~new_n560_ | ~\a[20] ) & (new_n560_ | \a[20] ))))) & (new_n561_ | (\a[17]  & ((new_n544_ ^ \a[20] ) | (new_n560_ & \a[20] ) | (~new_n67_ & (~new_n560_ | ~\a[20] ) & (new_n560_ | \a[20] ))) & ((new_n544_ & \a[20] ) | (~new_n544_ & ~\a[20] ) | ((~new_n560_ | ~\a[20] ) & (new_n67_ | (new_n560_ & \a[20] ) | (~new_n560_ & ~\a[20] ))))) | (~\a[17]  & ((new_n544_ ^ \a[20] ) ^ ((~new_n560_ | ~\a[20] ) & (new_n67_ | (new_n560_ & \a[20] ) | (~new_n560_ & ~\a[20] )))))));
endmodule


