// Benchmark "multiplier_675713_sat" written by ABC on Fri Jan 27 13:12:03 2023

module multiplier_675713_sat ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] ,
    \b[6] , \b[7] , \b[8] , \b[9] ,
    sat  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output sat;
  wire new_n33_, new_n34_, new_n35_, new_n36_, new_n37_, new_n38_, new_n39_,
    new_n40_, new_n41_, new_n42_, new_n43_, new_n44_, new_n45_, new_n46_,
    new_n47_, new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_,
    new_n54_, new_n55_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_,
    new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_,
    new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n74_,
    new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_,
    new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_,
    new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_,
    new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_;
  assign sat = ((~new_n257_ ^ new_n260_) | (new_n33_ & \a[2] ) | (~new_n221_ & (~new_n33_ | ~\a[2] ) & (new_n33_ | \a[2] ))) & ((~new_n257_ & new_n260_) | (new_n257_ & ~new_n260_) | ((~new_n33_ | ~\a[2] ) & (new_n221_ | (new_n33_ & \a[2] ) | (~new_n33_ & ~\a[2] )))) & ~new_n263_ & new_n264_ & (new_n221_ ^ (new_n33_ ^ \a[2] ));
  assign new_n33_ = ((~new_n34_ | ~\a[5] ) & ((new_n34_ & \a[5] ) | (~new_n34_ & ~\a[5] ) | ((~new_n161_ | ~\a[5] ) & (new_n171_ | (new_n161_ & \a[5] ) | (~new_n161_ & ~\a[5] ))))) ^ (~\a[5]  ^ (~new_n214_ ^ new_n220_));
  assign new_n34_ = ((\a[8]  & (((~new_n157_ | ~\a[11] ) & (((~new_n158_ | ~\a[11] ) & (new_n160_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] ))) | (new_n157_ & \a[11] ) | (~new_n157_ & ~\a[11] ))) | (new_n35_ & \a[11] ) | (~new_n35_ & ~\a[11] )) & ((new_n157_ & \a[11] ) | (((new_n158_ & \a[11] ) | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] ))) & (~new_n157_ | ~\a[11] ) & (new_n157_ | \a[11] )) | (new_n35_ ^ \a[11] ))) | (((\a[8]  & (((~new_n158_ | ~\a[11] ) & (new_n160_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] ))) | (new_n157_ & \a[11] ) | (~new_n157_ & ~\a[11] )) & ((new_n158_ & \a[11] ) | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] )) | (new_n157_ ^ \a[11] ))) | (((\a[8]  & (new_n160_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] )) & (~new_n160_ | (new_n158_ ^ \a[11] ))) | (~new_n95_ & (~\a[8]  | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] )) | (new_n160_ & (~new_n158_ ^ \a[11] ))) & (\a[8]  | (~new_n160_ ^ (new_n158_ ^ \a[11] ))))) & (~\a[8]  | (((new_n158_ & \a[11] ) | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] ))) & (~new_n157_ | ~\a[11] ) & (new_n157_ | \a[11] )) | ((~new_n158_ | ~\a[11] ) & (new_n160_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] )) & (~new_n157_ ^ \a[11] ))) & (\a[8]  | (((new_n158_ & \a[11] ) | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] ))) ^ (new_n157_ ^ \a[11] ))))) & (~\a[8]  | (((new_n157_ & \a[11] ) | (((new_n158_ & \a[11] ) | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] ))) & (~new_n157_ | ~\a[11] ) & (new_n157_ | \a[11] ))) & (~new_n35_ | ~\a[11] ) & (new_n35_ | \a[11] )) | ((~new_n157_ | ~\a[11] ) & (((~new_n158_ | ~\a[11] ) & (new_n160_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] ))) | (new_n157_ & \a[11] ) | (~new_n157_ & ~\a[11] )) & (~new_n35_ ^ \a[11] ))) & (\a[8]  | (((new_n157_ & \a[11] ) | (((new_n158_ & \a[11] ) | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] ))) & (~new_n157_ | ~\a[11] ) & (new_n157_ | \a[11] ))) ^ (new_n35_ ^ \a[11] ))))) ^ (\a[8]  ^ ((new_n152_ ^ \a[11] ) ^ ((new_n35_ & \a[11] ) | (((new_n157_ & \a[11] ) | (((new_n158_ & \a[11] ) | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] ))) & (~new_n157_ | ~\a[11] ) & (new_n157_ | \a[11] ))) & (~new_n35_ | ~\a[11] ) & (new_n35_ | \a[11] )))));
  assign new_n35_ = ~new_n70_ ^ (~new_n36_ ^ ~\a[14] );
  assign new_n36_ = new_n64_ ^ ((~new_n68_ & ~new_n69_) | (~new_n37_ & (new_n68_ | new_n69_) & (~new_n68_ | ~new_n69_)));
  assign new_n37_ = ~new_n38_ & ~new_n63_;
  assign new_n38_ = new_n59_ & (new_n39_ | (new_n58_ & (new_n43_ | (new_n57_ & (new_n46_ | (~new_n49_ & new_n56_))))));
  assign new_n39_ = (~\a[17]  ^ (new_n42_ & (~new_n40_ | ~new_n41_))) & ((\b[4]  & (~\a[17]  | ~\a[18] ) & (\a[17]  | \a[18] )) | (\b[3]  & \a[17]  & \a[18] ));
  assign new_n40_ = (\a[16]  | \a[17] ) & (~\a[16]  | ~\a[17] ) & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] );
  assign new_n41_ = ((\b[5]  & \b[6] ) | (((\b[4]  & \b[5] ) | (((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))) & (~\b[4]  | ~\b[5] ) & (\b[4]  | \b[5] ))) & (~\b[5]  | ~\b[6] ) & (\b[5]  | \b[6] ))) ^ (\b[6]  ^ \b[7] );
  assign new_n42_ = (~\b[5]  | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & (~\b[6]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[7]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ));
  assign new_n43_ = (~\a[17]  ^ (new_n45_ & (~new_n40_ | ~new_n44_))) & ((\b[3]  & (~\a[17]  | ~\a[18] ) & (\a[17]  | \a[18] )) | (\b[2]  & \a[17]  & \a[18] ));
  assign new_n44_ = ((\b[4]  & \b[5] ) | (((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))) & (~\b[4]  | ~\b[5] ) & (\b[4]  | \b[5] ))) ^ (\b[5]  ^ \b[6] );
  assign new_n45_ = (~\b[4]  | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & (~\b[5]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[6]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ));
  assign new_n46_ = (~\a[17]  ^ (new_n48_ & (~new_n40_ | ~new_n47_))) & ((\b[2]  & (~\a[17]  | ~\a[18] ) & (\a[17]  | \a[18] )) | (\b[1]  & \a[17]  & \a[18] ));
  assign new_n47_ = ((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))) ^ (\b[4]  ^ \b[5] );
  assign new_n48_ = (~\b[3]  | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & (~\b[4]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[5]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ));
  assign new_n49_ = (new_n52_ | (\a[17]  ^ (new_n51_ & (~new_n40_ | ~new_n50_)))) & ((~new_n53_ & (new_n54_ | ~new_n55_)) | (~new_n52_ & (~\a[17]  ^ (new_n51_ & (~new_n40_ | ~new_n50_)))) | (new_n52_ & (~\a[17]  | ~new_n51_ | (new_n40_ & new_n50_)) & (\a[17]  | (new_n51_ & (~new_n40_ | ~new_n50_)))));
  assign new_n50_ = (\b[3]  ^ \b[4] ) ^ ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] )));
  assign new_n51_ = (~\b[2]  | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & (~\b[3]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[4]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ));
  assign new_n52_ = (~\b[1]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[0]  | ~\a[17]  | ~\a[18] );
  assign new_n53_ = \b[0]  & (~\a[17]  | ~\a[18] ) & (\a[17]  | \a[18] ) & (~\b[0]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[1]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & ((~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\b[0]  ^ \b[1] )) & \a[17]  & (~\b[0]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[0]  | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & ((~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[1]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ));
  assign new_n54_ = \a[17]  ^ (((~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & (~\b[3]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[2]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )));
  assign new_n55_ = (\b[0]  & (~\a[17]  | ~\a[18] ) & (\a[17]  | \a[18] )) ^ ((~\b[0]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[1]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & ((~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\b[0]  ^ \b[1] )) & \a[17]  & (~\b[0]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[0]  | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & ((~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[1]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )));
  assign new_n56_ = (~\a[17]  ^ (new_n48_ & (~new_n40_ | ~new_n47_))) ^ ((\b[2]  & (~\a[17]  | ~\a[18] ) & (\a[17]  | \a[18] )) | (\b[1]  & \a[17]  & \a[18] ));
  assign new_n57_ = (~\a[17]  ^ (new_n45_ & (~new_n40_ | ~new_n44_))) ^ ((\b[3]  & (~\a[17]  | ~\a[18] ) & (\a[17]  | \a[18] )) | (\b[2]  & \a[17]  & \a[18] ));
  assign new_n58_ = (~\a[17]  ^ (new_n42_ & (~new_n40_ | ~new_n41_))) ^ ((\b[4]  & (~\a[17]  | ~\a[18] ) & (\a[17]  | \a[18] )) | (\b[3]  & \a[17]  & \a[18] ));
  assign new_n59_ = ~new_n62_ ^ (~\a[17]  ^ (new_n61_ & (~new_n40_ | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n60_ & (~\b[7]  ^ \b[8] )))));
  assign new_n60_ = (~\b[6]  | ~\b[7] ) & (((~\b[5]  | ~\b[6] ) & (((~\b[4]  | ~\b[5] ) & (((~\b[3]  | ~\b[4] ) & ((\b[3]  & \b[4] ) | (~\b[3]  & ~\b[4] ) | ((~\b[2]  | ~\b[3] ) & ((~\b[2]  & ~\b[3] ) | (\b[2]  & \b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] ))))) | (\b[4]  & \b[5] ) | (~\b[4]  & ~\b[5] ))) | (\b[5]  & \b[6] ) | (~\b[5]  & ~\b[6] ))) | (\b[6]  & \b[7] ) | (~\b[6]  & ~\b[7] ));
  assign new_n61_ = (~\b[6]  | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & (~\b[7]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[8]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ));
  assign new_n62_ = (~\b[5]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[4]  | ~\a[17]  | ~\a[18] );
  assign new_n63_ = ~new_n62_ & (~\a[17]  ^ (new_n61_ & (~new_n40_ | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n60_ & (~\b[7]  ^ \b[8] )))));
  assign new_n64_ = ~new_n65_ ^ ~new_n67_;
  assign new_n65_ = \a[17]  ^ (((new_n66_ ^ \b[9] ) | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[8]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[9]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )));
  assign new_n66_ = (~\b[8]  | ~\b[9] ) & ((~\b[8]  & ~\b[9] ) | (\b[8]  & \b[9] ) | ((~\b[7]  | ~\b[8] ) & (new_n60_ | (~\b[7]  & ~\b[8] ) | (\b[7]  & \b[8] ))));
  assign new_n67_ = (~\b[7]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[6]  | ~\a[17]  | ~\a[18] );
  assign new_n68_ = \a[17]  ^ (((\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n60_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[7]  | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[8]  | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[9]  | (\a[16]  ^ \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )));
  assign new_n69_ = (~\b[6]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[5]  | ~\a[17]  | ~\a[18] );
  assign new_n70_ = (~\a[14]  | (~new_n37_ & (~new_n68_ | ~new_n69_) & (new_n68_ | new_n69_)) | (new_n37_ & (~new_n68_ ^ new_n69_))) & (((new_n93_ | ~new_n94_) & (new_n71_ | (~new_n93_ & new_n94_) | (new_n93_ & ~new_n94_))) | (\a[14]  & (new_n37_ | (new_n68_ & new_n69_) | (~new_n68_ & ~new_n69_)) & (~new_n37_ | (new_n68_ ^ new_n69_))) | (~\a[14]  & (new_n37_ ^ (new_n68_ ^ new_n69_))));
  assign new_n71_ = (~new_n72_ | new_n91_) & (((~new_n73_ | new_n92_) & ((~new_n74_ & (new_n76_ | ~new_n90_)) | (new_n73_ & ~new_n92_) | (~new_n73_ & new_n92_))) | (new_n72_ & ~new_n91_) | (~new_n72_ & new_n91_));
  assign new_n72_ = new_n58_ ^ (new_n43_ | (new_n57_ & (new_n46_ | (~new_n49_ & new_n56_))));
  assign new_n73_ = new_n57_ ^ (new_n46_ | (~new_n49_ & new_n56_));
  assign new_n74_ = ~new_n75_ & (new_n49_ | ~new_n56_) & (~new_n49_ | new_n56_);
  assign new_n75_ = \a[14]  ^ (((\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n60_ & (~\b[7]  ^ \b[8] ))) & (~\b[7]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[8]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[6]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n76_ = (new_n77_ | ~new_n78_) & ((~new_n77_ & new_n78_) | (new_n77_ & ~new_n78_) | ((~new_n79_ | new_n80_) & ((~new_n79_ & new_n80_) | (new_n79_ & ~new_n80_) | ((new_n81_ | ~new_n89_) & (new_n82_ | (~new_n81_ & new_n89_) | (new_n81_ & ~new_n89_))))));
  assign new_n77_ = \a[14]  ^ ((~\b[6]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[7]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[5]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & (~new_n41_ | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )));
  assign new_n78_ = (new_n53_ | (~new_n54_ & new_n55_)) ^ (~new_n52_ ^ (~\a[17]  ^ (new_n51_ & (~new_n40_ | ~new_n50_))));
  assign new_n79_ = ~new_n54_ ^ new_n55_;
  assign new_n80_ = \a[14]  ^ ((~\b[5]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[6]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[4]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & (~new_n44_ | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )));
  assign new_n81_ = \a[14]  ^ ((~\b[4]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[5]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[3]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & (~new_n47_ | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )));
  assign new_n82_ = (~new_n85_ | (\a[14]  ^ (new_n84_ & (~new_n83_ | ~new_n50_)))) & ((~new_n86_ & (new_n87_ | ~new_n88_)) | (new_n85_ & (~\a[14]  ^ (new_n84_ & (~new_n83_ | ~new_n50_)))) | (~new_n85_ & (~\a[14]  | ~new_n84_ | (new_n83_ & new_n50_)) & (\a[14]  | (new_n84_ & (~new_n83_ | ~new_n50_)))));
  assign new_n83_ = (\a[13]  | \a[14] ) & (~\a[13]  | ~\a[14] ) & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] );
  assign new_n84_ = (~\b[3]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[4]  | (~\a[13]  ^ ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[2]  | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[12]  ^ ~\a[13] ));
  assign new_n85_ = ((\b[0]  & (\a[14]  ^ ~\a[15] ) & (\a[15]  | \a[16] ) & (~\a[15]  | ~\a[16] )) | (\b[1]  & (\a[16]  ^ ~\a[17] ) & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] )) | ((\a[16]  | \a[17] ) & (~\a[16]  | ~\a[17] ) & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ) & (\b[0]  ^ \b[1] ))) ^ (\a[17]  & \b[0]  & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] ));
  assign new_n86_ = \b[0]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] ) & (~\b[0]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[1]  | (~\a[13]  ^ ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\b[0]  ^ \b[1] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[13]  ^ ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[1]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[0]  | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[12]  ^ ~\a[13] ));
  assign new_n87_ = \a[14]  ^ (((~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[13]  ^ ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[2]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[1]  | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[12]  ^ ~\a[13] )));
  assign new_n88_ = (\b[0]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) ^ ((~\b[0]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[1]  | (~\a[13]  ^ ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\b[0]  ^ \b[1] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[13]  ^ ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[1]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[0]  | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[12]  ^ ~\a[13] )));
  assign new_n89_ = ((~\b[0]  | (~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  ^ ~\a[16] )) & (~\b[1]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[2]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & ((~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (\b[2]  ^ (\b[0]  | ~\b[1] )))) ^ (~\a[17]  | ((~\b[0]  | (~\a[14]  ^ ~\a[15] ) | (~\a[15]  & ~\a[16] ) | (\a[15]  & \a[16] )) & (~\b[1]  | (~\a[16]  ^ ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & ((~\a[16]  & ~\a[17] ) | (\a[16]  & \a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\b[0]  ^ \b[1] )) & \a[17]  & (~\b[0]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ))));
  assign new_n90_ = ~new_n75_ ^ (~new_n49_ ^ new_n56_);
  assign new_n91_ = \a[14]  ^ (((\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\b[9]  ^ ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))))))) & (~\b[8]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & (~\b[9]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )));
  assign new_n92_ = \a[14]  ^ (((\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n60_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[9]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[7]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )));
  assign new_n93_ = \a[14]  ^ (~\b[9]  | (((~\a[11]  ^ ~\a[12] ) | (~\a[12]  ^ ~\a[13] ) | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] )) & (new_n66_ | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ))));
  assign new_n94_ = new_n59_ ^ (new_n39_ | (new_n58_ & (new_n43_ | (new_n57_ & (new_n46_ | (~new_n49_ & new_n56_))))));
  assign new_n95_ = (~\a[8]  | (((new_n146_ & \a[11] ) | ((~new_n146_ | ~\a[11] ) & (new_n146_ | \a[11] ) & ((new_n147_ & ~new_n151_) | (~new_n148_ & (~new_n147_ | new_n151_) & (new_n147_ | ~new_n151_))))) & (~new_n144_ | ~\a[11] ) & (new_n144_ | \a[11] )) | ((~new_n146_ | ~\a[11] ) & ((new_n146_ & \a[11] ) | (~new_n146_ & ~\a[11] ) | ((~new_n147_ | new_n151_) & (new_n148_ | (new_n147_ & ~new_n151_) | (~new_n147_ & new_n151_)))) & (~new_n144_ ^ \a[11] ))) & (((~\a[8]  | ((~new_n146_ | ~\a[11] ) & (new_n146_ | \a[11] ) & ((new_n147_ & ~new_n151_) | (~new_n148_ & (~new_n147_ | new_n151_) & (new_n147_ | ~new_n151_)))) | ((~new_n146_ ^ \a[11] ) & (~new_n147_ | new_n151_) & (new_n148_ | (new_n147_ & ~new_n151_) | (~new_n147_ & new_n151_)))) & (((~\a[8]  | (~new_n148_ & (~new_n147_ | new_n151_) & (new_n147_ | ~new_n151_)) | (new_n148_ & (~new_n147_ ^ ~new_n151_))) & (new_n96_ | (\a[8]  & (new_n148_ | (new_n147_ & ~new_n151_) | (~new_n147_ & new_n151_)) & (~new_n148_ | (new_n147_ ^ ~new_n151_))) | (~\a[8]  & (new_n148_ ^ (new_n147_ ^ ~new_n151_))))) | (\a[8]  & ((new_n146_ & \a[11] ) | (~new_n146_ & ~\a[11] ) | ((~new_n147_ | new_n151_) & (new_n148_ | (new_n147_ & ~new_n151_) | (~new_n147_ & new_n151_)))) & ((new_n146_ ^ \a[11] ) | (new_n147_ & ~new_n151_) | (~new_n148_ & (~new_n147_ | new_n151_) & (new_n147_ | ~new_n151_)))) | (~\a[8]  & ((~new_n146_ ^ \a[11] ) ^ ((new_n147_ & ~new_n151_) | (~new_n148_ & (~new_n147_ | new_n151_) & (new_n147_ | ~new_n151_))))))) | (\a[8]  & (((~new_n146_ | ~\a[11] ) & ((new_n146_ & \a[11] ) | (~new_n146_ & ~\a[11] ) | ((~new_n147_ | new_n151_) & (new_n148_ | (new_n147_ & ~new_n151_) | (~new_n147_ & new_n151_))))) | (new_n144_ & \a[11] ) | (~new_n144_ & ~\a[11] )) & ((new_n146_ & \a[11] ) | ((~new_n146_ | ~\a[11] ) & (new_n146_ | \a[11] ) & ((new_n147_ & ~new_n151_) | (~new_n148_ & (~new_n147_ | new_n151_) & (new_n147_ | ~new_n151_)))) | (new_n144_ ^ \a[11] ))) | (~\a[8]  & (((~new_n146_ | ~\a[11] ) & ((new_n146_ & \a[11] ) | (~new_n146_ & ~\a[11] ) | ((~new_n147_ | new_n151_) & (new_n148_ | (new_n147_ & ~new_n151_) | (~new_n147_ & new_n151_))))) ^ (new_n144_ ^ \a[11] ))));
  assign new_n96_ = (~new_n97_ | ~\a[8] ) & ((new_n97_ & \a[8] ) | (~new_n97_ & ~\a[8] ) | ((~new_n118_ | ~\a[8] ) & ((new_n118_ & \a[8] ) | (~new_n118_ & ~\a[8] ) | (~new_n119_ & (new_n121_ | ~new_n143_)))));
  assign new_n97_ = new_n115_ ^ (new_n98_ | (~new_n98_ & ~new_n114_ & ((~new_n117_ & (new_n82_ | (~new_n81_ & new_n89_) | (new_n81_ & ~new_n89_)) & (~new_n82_ | (~new_n81_ ^ new_n89_))) | (~new_n100_ & (new_n117_ | (~new_n82_ & (new_n81_ | ~new_n89_) & (~new_n81_ | new_n89_)) | (new_n82_ & (new_n81_ ^ new_n89_))) & (~new_n117_ | (~new_n82_ ^ (~new_n81_ ^ new_n89_)))))));
  assign new_n98_ = ~new_n99_ & ((~new_n79_ & new_n80_) | (new_n79_ & ~new_n80_) | ((new_n81_ | ~new_n89_) & (new_n82_ | (~new_n81_ & new_n89_) | (new_n81_ & ~new_n89_)))) & ((~new_n79_ ^ new_n80_) | (~new_n81_ & new_n89_) | (~new_n82_ & (new_n81_ | ~new_n89_) & (~new_n81_ | new_n89_)));
  assign new_n99_ = \a[11]  ^ (((\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n60_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[9]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[7]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n100_ = (new_n101_ | ~new_n102_) & ((~new_n101_ & new_n102_) | (new_n101_ & ~new_n102_) | ((~new_n103_ | new_n104_) & ((~new_n103_ & new_n104_) | (new_n103_ & ~new_n104_) | ((new_n105_ | ~new_n113_) & (new_n106_ | (~new_n105_ & new_n113_) | (new_n105_ & ~new_n113_))))));
  assign new_n101_ = \a[11]  ^ ((~new_n41_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[6]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[7]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[5]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n102_ = (new_n86_ | (~new_n87_ & new_n88_)) ^ (new_n85_ ^ (~\a[14]  ^ (new_n84_ & (~new_n83_ | ~new_n50_))));
  assign new_n103_ = ~new_n87_ ^ new_n88_;
  assign new_n104_ = \a[11]  ^ ((~new_n44_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[5]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[6]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[4]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n105_ = \a[11]  ^ ((~new_n47_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[4]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[5]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[3]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n106_ = (~new_n109_ | (\a[11]  ^ (new_n108_ & (~new_n50_ | ~new_n107_)))) & ((~new_n110_ & (new_n111_ | ~new_n112_)) | (new_n109_ & (~\a[11]  ^ (new_n108_ & (~new_n50_ | ~new_n107_)))) | (~new_n109_ & (~\a[11]  | ~new_n108_ | (new_n50_ & new_n107_)) & (\a[11]  | (new_n108_ & (~new_n50_ | ~new_n107_)))));
  assign new_n107_ = (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] ) & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] );
  assign new_n108_ = (~\b[3]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[4]  | (~\a[10]  ^ ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[2]  | (~\a[9]  ^ ~\a[10] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] ));
  assign new_n109_ = ((\b[0]  & (\a[11]  ^ ~\a[12] ) & (\a[12]  | \a[13] ) & (~\a[12]  | ~\a[13] )) | (\b[1]  & (\a[13]  ^ ~\a[14] ) & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] )) | ((\a[13]  | \a[14] ) & (~\a[13]  | ~\a[14] ) & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ) & (\b[0]  ^ \b[1] ))) ^ (\a[14]  & \b[0]  & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ));
  assign new_n110_ = \b[0]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] ) & (~\b[0]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (~\a[10]  ^ ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\b[0]  ^ \b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[10]  ^ ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[1]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[0]  | (~\a[9]  ^ ~\a[10] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] ));
  assign new_n111_ = \a[11]  ^ (((~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[10]  ^ ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[2]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (~\a[9]  ^ ~\a[10] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n112_ = (\b[0]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] )) ^ ((~\b[0]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (~\a[10]  ^ ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\b[0]  ^ \b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[10]  ^ ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[1]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[0]  | (~\a[9]  ^ ~\a[10] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n113_ = (~\a[14]  | ((~\b[0]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[1]  | (~\a[13]  ^ ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\b[0]  ^ \b[1] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )))) ^ ((~\b[0]  | (~\a[11]  ^ ~\a[12] ) | (~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[12]  ^ ~\a[13] )) & (~\b[1]  | (~\a[11]  ^ ~\a[12] ) | (~\a[12]  & ~\a[13] ) | (\a[12]  & \a[13] )) & (~\b[2]  | (~\a[13]  ^ ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((~\a[13]  & ~\a[14] ) | (\a[13]  & \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))));
  assign new_n114_ = new_n99_ & ((new_n79_ ^ new_n80_) ^ ((~new_n81_ & new_n89_) | (~new_n82_ & (new_n81_ | ~new_n89_) & (~new_n81_ | new_n89_))));
  assign new_n115_ = ~new_n116_ ^ ((~new_n77_ ^ new_n78_) ^ ((new_n79_ & ~new_n80_) | ((new_n79_ | ~new_n80_) & (~new_n79_ | new_n80_) & ((~new_n81_ & new_n89_) | (~new_n82_ & (new_n81_ | ~new_n89_) & (~new_n81_ | new_n89_))))));
  assign new_n116_ = \a[11]  ^ (((\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\b[9]  ^ ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))))))) & (~\b[9]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[8]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n117_ = \a[11]  ^ (((\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n60_ & (~\b[7]  ^ \b[8] ))) & (~\b[7]  | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[8]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[6]  | (~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n118_ = (~new_n98_ & ~new_n114_) ^ ((~new_n117_ & (new_n82_ | (~new_n81_ & new_n89_) | (new_n81_ & ~new_n89_)) & (~new_n82_ | (~new_n81_ ^ new_n89_))) | (~new_n100_ & (new_n117_ | (~new_n82_ & (new_n81_ | ~new_n89_) & (~new_n81_ | new_n89_)) | (new_n82_ & (new_n81_ ^ new_n89_))) & (~new_n117_ | (~new_n82_ ^ (~new_n81_ ^ new_n89_)))));
  assign new_n119_ = (new_n100_ | ~new_n120_) & (~new_n100_ | new_n120_) & (~\a[8]  ^ (~\b[9]  | ((new_n66_ | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & ((\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )))));
  assign new_n120_ = ~new_n117_ ^ (~new_n82_ ^ (~new_n81_ ^ new_n89_));
  assign new_n121_ = (~new_n123_ | new_n141_) & ((new_n123_ & ~new_n141_) | (~new_n123_ & new_n141_) | (~new_n124_ & (((new_n142_ | (new_n122_ & ~new_n106_) | (~new_n122_ & new_n106_)) & (new_n126_ | (~new_n142_ & (~new_n122_ | new_n106_) & (new_n122_ | ~new_n106_)) | (new_n142_ & (~new_n122_ ^ ~new_n106_)))) | new_n124_ | new_n140_)));
  assign new_n122_ = ~new_n105_ ^ new_n113_;
  assign new_n123_ = (~new_n101_ ^ new_n102_) ^ ((new_n103_ & ~new_n104_) | ((new_n103_ | ~new_n104_) & (~new_n103_ | new_n104_) & ((~new_n105_ & new_n113_) | (~new_n106_ & (new_n105_ | ~new_n113_) & (~new_n105_ | new_n113_)))));
  assign new_n124_ = ~new_n125_ & ((~new_n103_ & new_n104_) | (new_n103_ & ~new_n104_) | ((new_n105_ | ~new_n113_) & (new_n106_ | (~new_n105_ & new_n113_) | (new_n105_ & ~new_n113_)))) & ((~new_n103_ ^ new_n104_) | (~new_n105_ & new_n113_) | (~new_n106_ & (new_n105_ | ~new_n113_) & (~new_n105_ | new_n113_)));
  assign new_n125_ = \a[8]  ^ (((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n60_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[9]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[7]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n126_ = (~new_n127_ | new_n128_) & ((~new_n127_ & new_n128_) | (new_n127_ & ~new_n128_) | ((~new_n129_ | new_n130_) & ((~new_n129_ & new_n130_) | (new_n129_ & ~new_n130_) | ((new_n131_ | ~new_n139_) & (new_n132_ | (~new_n131_ & new_n139_) | (new_n131_ & ~new_n139_))))));
  assign new_n127_ = (new_n110_ | (~new_n111_ & new_n112_)) ^ (new_n109_ ^ (~\a[11]  ^ (new_n108_ & (~new_n50_ | ~new_n107_))));
  assign new_n128_ = \a[8]  ^ ((~new_n41_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[6]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[7]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[5]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n129_ = ~new_n111_ ^ new_n112_;
  assign new_n130_ = \a[8]  ^ ((~new_n44_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[5]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[6]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[4]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n131_ = \a[8]  ^ ((~new_n47_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[4]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[5]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[3]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n132_ = (~new_n135_ | (\a[8]  ^ (new_n134_ & (~new_n50_ | ~new_n133_)))) & ((~new_n136_ & (new_n137_ | ~new_n138_)) | (new_n135_ & (~\a[8]  ^ (new_n134_ & (~new_n50_ | ~new_n133_)))) | (~new_n135_ & (~\a[8]  | ~new_n134_ | (new_n50_ & new_n133_)) & (\a[8]  | (new_n134_ & (~new_n50_ | ~new_n133_)))));
  assign new_n133_ = (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] ) & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] );
  assign new_n134_ = (~\b[3]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[4]  | (~\a[7]  ^ ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[2]  | (~\a[6]  ^ ~\a[7] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  ^ ~\a[6] ));
  assign new_n135_ = ((\b[0]  & (\a[8]  ^ ~\a[9] ) & (\a[9]  | \a[10] ) & (~\a[9]  | ~\a[10] )) | (\b[1]  & (\a[10]  ^ ~\a[11] ) & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] )) | ((\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] ) & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\b[0]  ^ \b[1] ))) ^ (\a[11]  & \b[0]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ));
  assign new_n136_ = \b[0]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] ) & (~\b[0]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[7]  ^ ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\b[0]  ^ \b[1] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[7]  ^ ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[1]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  ^ ~\a[6] ));
  assign new_n137_ = \a[8]  ^ (((~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[7]  ^ ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[2]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[6]  ^ ~\a[7] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n138_ = (\b[0]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] )) ^ ((~\b[0]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[7]  ^ ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\b[0]  ^ \b[1] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[7]  ^ ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[1]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n139_ = (~\a[11]  | ((~\b[0]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (~\a[10]  ^ ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\b[0]  ^ \b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )))) ^ ((~\b[1]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[2]  | (~\a[10]  ^ ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[9]  ^ ~\a[10] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n140_ = new_n125_ & ((new_n103_ ^ new_n104_) ^ ((~new_n105_ & new_n113_) | (~new_n106_ & (new_n105_ | ~new_n113_) & (~new_n105_ | new_n113_))));
  assign new_n141_ = \a[8]  ^ (((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\b[9]  ^ ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))))))) & (~\b[9]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[8]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n142_ = \a[8]  ^ (((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n60_ & (~\b[7]  ^ \b[8] ))) & (~\b[7]  | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[8]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[6]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n143_ = (~new_n100_ ^ new_n120_) ^ (~\a[8]  ^ (~\b[9]  | ((new_n66_ | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )) & ((\a[6]  ^ \a[7] ) | (\a[5]  ^ \a[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] )))));
  assign new_n144_ = new_n145_ ^ ((new_n73_ & ~new_n92_) | ((~new_n73_ | new_n92_) & (new_n73_ | ~new_n92_) & (new_n74_ | (~new_n76_ & new_n90_))));
  assign new_n145_ = ~new_n91_ ^ (new_n58_ ^ (new_n43_ | (new_n57_ & (new_n46_ | (~new_n49_ & new_n56_)))));
  assign new_n146_ = (new_n74_ | (~new_n76_ & new_n90_)) ^ (new_n73_ ^ ~new_n92_);
  assign new_n147_ = ~new_n76_ ^ new_n90_;
  assign new_n148_ = (~new_n150_ | new_n116_) & ((new_n150_ & ~new_n116_) | (~new_n150_ & new_n116_) | (~new_n98_ & (((new_n117_ | (new_n149_ & ~new_n82_) | (~new_n149_ & new_n82_)) & (new_n100_ | (~new_n117_ & (~new_n149_ | new_n82_) & (new_n149_ | ~new_n82_)) | (new_n117_ & (~new_n149_ ^ ~new_n82_)))) | new_n98_ | new_n114_)));
  assign new_n149_ = ~new_n81_ ^ new_n89_;
  assign new_n150_ = (~new_n77_ ^ new_n78_) ^ ((new_n79_ & ~new_n80_) | ((new_n79_ | ~new_n80_) & (~new_n79_ | new_n80_) & ((~new_n81_ & new_n89_) | (~new_n82_ & (new_n81_ | ~new_n89_) & (~new_n81_ | new_n89_)))));
  assign new_n151_ = \a[11]  ^ (~\b[9]  | ((new_n66_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((~\a[9]  ^ ~\a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] ))));
  assign new_n152_ = ((new_n36_ & \a[14] ) | (~new_n70_ & (~new_n36_ | ~\a[14] ) & (new_n36_ | \a[14] ))) ^ (\a[14]  ^ (~new_n153_ ^ new_n154_));
  assign new_n153_ = (new_n65_ | new_n67_) & (((new_n68_ | new_n69_) & (new_n37_ | (~new_n68_ & ~new_n69_) | (new_n68_ & new_n69_))) | (~new_n65_ & ~new_n67_) | (new_n65_ & new_n67_));
  assign new_n154_ = ~new_n155_ ^ ~new_n156_;
  assign new_n155_ = \a[17]  ^ (~\b[9]  | (((\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[15]  ^ ~\a[16] ) | (~\a[14]  ^ ~\a[15] )) & (new_n66_ | (\a[16]  & \a[17] ) | (~\a[16]  & ~\a[17] ) | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ))));
  assign new_n156_ = (~\b[8]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )) & (~\b[7]  | ~\a[17]  | ~\a[18] );
  assign new_n157_ = ((~new_n93_ & new_n94_) | (~new_n71_ & (new_n93_ | ~new_n94_) & (~new_n93_ | new_n94_))) ^ (\a[14]  ^ (~new_n37_ ^ (new_n68_ ^ new_n69_)));
  assign new_n158_ = ~new_n71_ ^ new_n159_;
  assign new_n159_ = ~new_n93_ ^ new_n94_;
  assign new_n160_ = (~new_n144_ | ~\a[11] ) & ((new_n144_ & \a[11] ) | (~new_n144_ & ~\a[11] ) | ((~new_n146_ | ~\a[11] ) & ((new_n146_ & \a[11] ) | (~new_n146_ & ~\a[11] ) | ((~new_n147_ | new_n151_) & (new_n148_ | (new_n147_ & ~new_n151_) | (~new_n147_ & new_n151_))))));
  assign new_n161_ = new_n170_ ^ (new_n162_ | (~new_n165_ & new_n169_));
  assign new_n162_ = \a[8]  & (new_n163_ | ~new_n164_) & (~new_n163_ | new_n164_);
  assign new_n163_ = (~\a[11]  | (~new_n71_ & new_n159_) | (new_n71_ & ~new_n159_)) & (((~new_n144_ | ~\a[11] ) & ((new_n144_ & \a[11] ) | (~new_n144_ & ~\a[11] ) | ((~new_n146_ | ~\a[11] ) & ((new_n146_ & \a[11] ) | (~new_n146_ & ~\a[11] ) | ((~new_n147_ | new_n151_) & (new_n148_ | (~new_n147_ & new_n151_) | (new_n147_ & ~new_n151_))))))) | (\a[11]  & (new_n71_ | ~new_n159_) & (~new_n71_ | new_n159_)) | (~\a[11]  & (new_n71_ ^ new_n159_)));
  assign new_n164_ = \a[11]  ^ (((~new_n93_ & new_n94_) | (~new_n71_ & (new_n93_ | ~new_n94_) & (~new_n93_ | new_n94_))) ^ (\a[14]  ^ (~new_n37_ ^ (new_n68_ ^ new_n69_))));
  assign new_n165_ = (~new_n166_ | ~\a[8] ) & ((new_n166_ & \a[8] ) | (~new_n166_ & ~\a[8] ) | ((~new_n167_ | ~\a[8] ) & ((new_n167_ & \a[8] ) | (~new_n167_ & ~\a[8] ) | ((~\a[8]  | (new_n168_ & ((new_n147_ & ~new_n151_) | (~new_n148_ & (new_n147_ | ~new_n151_) & (~new_n147_ | new_n151_)))) | (~new_n168_ & (~new_n147_ | new_n151_) & (new_n148_ | (~new_n147_ & new_n151_) | (new_n147_ & ~new_n151_)))) & (((~\a[8]  | (~new_n148_ & (new_n147_ | ~new_n151_) & (~new_n147_ | new_n151_)) | (new_n148_ & (new_n147_ ^ new_n151_))) & (new_n96_ | (\a[8]  & (new_n148_ | (~new_n147_ & new_n151_) | (new_n147_ & ~new_n151_)) & (~new_n148_ | (~new_n147_ ^ new_n151_))) | (~\a[8]  & (new_n148_ ^ (~new_n147_ ^ new_n151_))))) | (\a[8]  & (~new_n168_ | ((~new_n147_ | new_n151_) & (new_n148_ | (~new_n147_ & new_n151_) | (new_n147_ & ~new_n151_)))) & (new_n168_ | (new_n147_ & ~new_n151_) | (~new_n148_ & (new_n147_ | ~new_n151_) & (~new_n147_ | new_n151_)))) | (~\a[8]  & (~new_n168_ ^ ((new_n147_ & ~new_n151_) | (~new_n148_ & (new_n147_ | ~new_n151_) & (~new_n147_ | new_n151_))))))))));
  assign new_n166_ = ((new_n144_ & \a[11] ) | ((~new_n144_ | ~\a[11] ) & (new_n144_ | \a[11] ) & ((new_n146_ & \a[11] ) | ((~new_n146_ | ~\a[11] ) & (new_n146_ | \a[11] ) & ((new_n147_ & ~new_n151_) | (~new_n148_ & (new_n147_ | ~new_n151_) & (~new_n147_ | new_n151_))))))) ^ (\a[11]  ^ (~new_n71_ ^ new_n159_));
  assign new_n167_ = (new_n144_ ^ \a[11] ) ^ ((new_n146_ & \a[11] ) | ((~new_n146_ | ~\a[11] ) & (new_n146_ | \a[11] ) & ((new_n147_ & ~new_n151_) | (~new_n148_ & (~new_n147_ | new_n151_) & (new_n147_ | ~new_n151_)))));
  assign new_n168_ = \a[11]  ^ ((new_n74_ | (~new_n76_ & new_n90_)) ^ (new_n73_ ^ ~new_n92_));
  assign new_n169_ = \a[8]  ^ (~new_n163_ ^ new_n164_);
  assign new_n170_ = \a[8]  ^ (((new_n157_ & \a[11] ) | (~new_n163_ & (~new_n157_ | ~\a[11] ) & (new_n157_ | \a[11] ))) ^ (\a[11]  ^ (~new_n70_ ^ (new_n36_ ^ \a[14] ))));
  assign new_n171_ = (~\a[5]  | (~new_n165_ & new_n169_) | (new_n165_ & ~new_n169_)) & (((~new_n172_ | ~\a[5] ) & (((~new_n173_ | ~\a[5] ) & (new_n174_ | (new_n173_ & \a[5] ) | (~new_n173_ & ~\a[5] ))) | (new_n172_ & \a[5] ) | (~new_n172_ & ~\a[5] ))) | (\a[5]  & (new_n165_ | ~new_n169_) & (~new_n165_ | new_n169_)) | (~\a[5]  & (new_n165_ ^ new_n169_)));
  assign new_n172_ = (new_n166_ ^ \a[8] ) ^ ((new_n167_ & \a[8] ) | ((~new_n167_ | ~\a[8] ) & (new_n167_ | \a[8] ) & ((\a[8]  & (~new_n168_ | ((~new_n147_ | new_n151_) & (new_n148_ | (~new_n147_ & new_n151_) | (new_n147_ & ~new_n151_)))) & (new_n168_ | (new_n147_ & ~new_n151_) | (~new_n148_ & (new_n147_ | ~new_n151_) & (~new_n147_ | new_n151_)))) | (((\a[8]  & (new_n148_ | (~new_n147_ & new_n151_) | (new_n147_ & ~new_n151_)) & (~new_n148_ | (~new_n147_ ^ new_n151_))) | (~new_n96_ & (~\a[8]  | (~new_n148_ & (new_n147_ | ~new_n151_) & (~new_n147_ | new_n151_)) | (new_n148_ & (new_n147_ ^ new_n151_))) & (\a[8]  | (~new_n148_ ^ (~new_n147_ ^ new_n151_))))) & (~\a[8]  | (new_n168_ & ((new_n147_ & ~new_n151_) | (~new_n148_ & (new_n147_ | ~new_n151_) & (~new_n147_ | new_n151_)))) | (~new_n168_ & (~new_n147_ | new_n151_) & (new_n148_ | (~new_n147_ & new_n151_) | (new_n147_ & ~new_n151_)))) & (\a[8]  | (new_n168_ ^ ((new_n147_ & ~new_n151_) | (~new_n148_ & (new_n147_ | ~new_n151_) & (~new_n147_ | new_n151_)))))))));
  assign new_n173_ = ((\a[8]  & ((new_n146_ & \a[11] ) | (~new_n146_ & ~\a[11] ) | ((~new_n147_ | new_n151_) & (new_n148_ | (new_n147_ & ~new_n151_) | (~new_n147_ & new_n151_)))) & ((new_n146_ ^ \a[11] ) | (new_n147_ & ~new_n151_) | (~new_n148_ & (~new_n147_ | new_n151_) & (new_n147_ | ~new_n151_)))) | (((\a[8]  & (new_n148_ | (new_n147_ & ~new_n151_) | (~new_n147_ & new_n151_)) & (~new_n148_ | (new_n147_ ^ ~new_n151_))) | (~new_n96_ & (~\a[8]  | (~new_n148_ & (~new_n147_ | new_n151_) & (new_n147_ | ~new_n151_)) | (new_n148_ & (~new_n147_ ^ ~new_n151_))) & (\a[8]  | (~new_n148_ ^ (new_n147_ ^ ~new_n151_))))) & (~\a[8]  | ((~new_n146_ | ~\a[11] ) & (new_n146_ | \a[11] ) & ((new_n147_ & ~new_n151_) | (~new_n148_ & (~new_n147_ | new_n151_) & (new_n147_ | ~new_n151_)))) | ((~new_n146_ ^ \a[11] ) & (~new_n147_ | new_n151_) & (new_n148_ | (new_n147_ & ~new_n151_) | (~new_n147_ & new_n151_)))) & (\a[8]  | ((new_n146_ ^ \a[11] ) ^ ((new_n147_ & ~new_n151_) | (~new_n148_ & (~new_n147_ | new_n151_) & (new_n147_ | ~new_n151_))))))) ^ (\a[8]  ^ (((new_n146_ & \a[11] ) | ((~new_n146_ | ~\a[11] ) & (new_n146_ | \a[11] ) & ((new_n147_ & ~new_n151_) | (~new_n148_ & (~new_n147_ | new_n151_) & (new_n147_ | ~new_n151_))))) ^ (new_n144_ ^ \a[11] )));
  assign new_n174_ = (~\a[5]  | (~new_n175_ & new_n177_) | (new_n175_ & ~new_n177_)) & ((\a[5]  & (new_n175_ | ~new_n177_) & (~new_n175_ | new_n177_)) | (~\a[5]  & (new_n175_ ^ new_n177_)) | ((~new_n178_ | ~\a[5] ) & ((new_n178_ & \a[5] ) | (~new_n178_ & ~\a[5] ) | ((~new_n179_ | ~\a[5] ) & ((new_n179_ & \a[5] ) | (~new_n179_ & ~\a[5] ) | (~new_n180_ & (new_n181_ | ~new_n213_)))))));
  assign new_n175_ = (~\a[8]  | (~new_n148_ & new_n176_) | (new_n148_ & ~new_n176_)) & ((\a[8]  & (new_n148_ | ~new_n176_) & (~new_n148_ | new_n176_)) | (~\a[8]  & (new_n148_ ^ new_n176_)) | ((~new_n97_ | ~\a[8] ) & ((new_n97_ & \a[8] ) | (~new_n97_ & ~\a[8] ) | ((~new_n118_ | ~\a[8] ) & ((new_n118_ & \a[8] ) | (~new_n118_ & ~\a[8] ) | (~new_n119_ & (new_n121_ | ~new_n143_)))))));
  assign new_n176_ = ~new_n151_ ^ (~new_n76_ ^ new_n90_);
  assign new_n177_ = \a[8]  ^ (new_n168_ ^ ((new_n147_ & ~new_n151_) | (~new_n148_ & (new_n147_ | ~new_n151_) & (~new_n147_ | new_n151_))));
  assign new_n178_ = (\a[8]  ^ (~new_n148_ ^ new_n176_)) ^ ((new_n97_ & \a[8] ) | ((~new_n97_ | ~\a[8] ) & (new_n97_ | \a[8] ) & ((new_n118_ & \a[8] ) | ((~new_n118_ | ~\a[8] ) & (new_n118_ | \a[8] ) & (new_n119_ | (~new_n121_ & new_n143_))))));
  assign new_n179_ = (new_n97_ ^ \a[8] ) ^ ((new_n118_ & \a[8] ) | ((~new_n118_ | ~\a[8] ) & (new_n118_ | \a[8] ) & (new_n119_ | (~new_n121_ & new_n143_))));
  assign new_n180_ = \a[5]  & ((new_n118_ & \a[8] ) | (~new_n118_ & ~\a[8] ) | (~new_n119_ & (new_n121_ | ~new_n143_))) & ((new_n118_ ^ \a[8] ) | new_n119_ | (~new_n121_ & new_n143_));
  assign new_n181_ = (~\a[5]  | (~new_n121_ & new_n143_) | (new_n121_ & ~new_n143_)) & ((\a[5]  & (new_n121_ | ~new_n143_) & (~new_n121_ | new_n143_)) | (~\a[5]  & (new_n121_ ^ new_n143_)) | ((~new_n182_ | ~\a[5] ) & ((new_n182_ & \a[5] ) | (~new_n182_ & ~\a[5] ) | ((~new_n185_ | ~\a[5] ) & ((new_n185_ & \a[5] ) | (~new_n185_ & ~\a[5] ) | (~new_n186_ & (new_n189_ | ~new_n212_)))))));
  assign new_n182_ = new_n184_ ^ ((~new_n125_ & (~new_n183_ | ((new_n105_ | ~new_n113_) & (new_n106_ | (~new_n105_ & new_n113_) | (new_n105_ & ~new_n113_)))) & (new_n183_ | (~new_n105_ & new_n113_) | (~new_n106_ & (new_n105_ | ~new_n113_) & (~new_n105_ | new_n113_)))) | (((~new_n142_ & (new_n106_ | (~new_n105_ & new_n113_) | (new_n105_ & ~new_n113_)) & (~new_n106_ | (~new_n105_ ^ new_n113_))) | (~new_n126_ & (new_n142_ | (~new_n106_ & (new_n105_ | ~new_n113_) & (~new_n105_ | new_n113_)) | (new_n106_ & (new_n105_ ^ new_n113_))) & (~new_n142_ | (~new_n106_ ^ (~new_n105_ ^ new_n113_))))) & (new_n125_ | (new_n183_ & ((~new_n105_ & new_n113_) | (~new_n106_ & (new_n105_ | ~new_n113_) & (~new_n105_ | new_n113_)))) | (~new_n183_ & (new_n105_ | ~new_n113_) & (new_n106_ | (~new_n105_ & new_n113_) | (new_n105_ & ~new_n113_)))) & (~new_n125_ | (new_n183_ ^ ((~new_n105_ & new_n113_) | (~new_n106_ & (new_n105_ | ~new_n113_) & (~new_n105_ | new_n113_)))))));
  assign new_n183_ = ~new_n103_ ^ new_n104_;
  assign new_n184_ = ~new_n141_ ^ ((~new_n101_ ^ new_n102_) ^ ((new_n103_ & ~new_n104_) | ((new_n103_ | ~new_n104_) & (~new_n103_ | new_n104_) & ((~new_n105_ & new_n113_) | (~new_n106_ & (new_n105_ | ~new_n113_) & (~new_n105_ | new_n113_))))));
  assign new_n185_ = (~new_n124_ & ~new_n140_) ^ ((~new_n142_ & (new_n106_ | (~new_n105_ & new_n113_) | (new_n105_ & ~new_n113_)) & (~new_n106_ | (~new_n105_ ^ new_n113_))) | (~new_n126_ & (new_n142_ | (~new_n106_ & (new_n105_ | ~new_n113_) & (~new_n105_ | new_n113_)) | (new_n106_ & (new_n105_ ^ new_n113_))) & (~new_n142_ | (~new_n106_ ^ (~new_n105_ ^ new_n113_)))));
  assign new_n186_ = ~new_n188_ & (new_n126_ | ~new_n187_) & (~new_n126_ | new_n187_);
  assign new_n187_ = ~new_n142_ ^ (~new_n106_ ^ (~new_n105_ ^ new_n113_));
  assign new_n188_ = \a[5]  ^ (~\b[9]  | ((new_n66_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] ))));
  assign new_n189_ = (~new_n191_ | new_n210_) & ((new_n191_ & ~new_n210_) | (~new_n191_ & new_n210_) | (~new_n192_ & (new_n192_ | new_n194_ | ((new_n211_ | (new_n190_ & ~new_n132_) | (~new_n190_ & new_n132_)) & (new_n195_ | (~new_n211_ & (~new_n190_ | new_n132_) & (new_n190_ | ~new_n132_)) | (new_n211_ & (~new_n190_ ^ ~new_n132_)))))));
  assign new_n190_ = ~new_n131_ ^ new_n139_;
  assign new_n191_ = (~new_n127_ ^ new_n128_) ^ ((new_n129_ & ~new_n130_) | ((new_n129_ | ~new_n130_) & (~new_n129_ | new_n130_) & ((~new_n131_ & new_n139_) | (~new_n132_ & (new_n131_ | ~new_n139_) & (~new_n131_ | new_n139_)))));
  assign new_n192_ = ~new_n193_ & ((~new_n129_ & new_n130_) | (new_n129_ & ~new_n130_) | ((new_n131_ | ~new_n139_) & (new_n132_ | (~new_n131_ & new_n139_) | (new_n131_ & ~new_n139_)))) & ((~new_n129_ ^ new_n130_) | (~new_n131_ & new_n139_) | (~new_n132_ & (new_n131_ | ~new_n139_) & (~new_n131_ | new_n139_)));
  assign new_n193_ = \a[5]  ^ (((\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n60_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[8]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[9]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[7]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n194_ = new_n193_ & ((new_n129_ ^ new_n130_) ^ ((~new_n131_ & new_n139_) | (~new_n132_ & (new_n131_ | ~new_n139_) & (~new_n131_ | new_n139_))));
  assign new_n195_ = (~new_n196_ | new_n197_) & ((~new_n196_ & new_n197_) | (new_n196_ & ~new_n197_) | ((~new_n198_ | new_n199_) & ((~new_n198_ & new_n199_) | (new_n198_ & ~new_n199_) | ((new_n200_ | ~new_n209_) & (new_n203_ | (~new_n200_ & new_n209_) | (new_n200_ & ~new_n209_))))));
  assign new_n196_ = (new_n136_ | (~new_n137_ & new_n138_)) ^ (new_n135_ ^ (~\a[8]  ^ (new_n134_ & (~new_n50_ | ~new_n133_))));
  assign new_n197_ = \a[5]  ^ ((~new_n41_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[6]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[7]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[5]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n198_ = ~new_n137_ ^ new_n138_;
  assign new_n199_ = \a[5]  ^ ((~new_n44_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[5]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[6]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[4]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n200_ = \a[5]  ^ (new_n202_ & (~new_n47_ | ~new_n201_));
  assign new_n201_ = (\a[4]  | \a[5] ) & (~\a[4]  | ~\a[5] ) & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] );
  assign new_n202_ = (~\b[4]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[5]  | (~\a[4]  ^ ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[3]  | (~\a[3]  ^ ~\a[4] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  ^ ~\a[3] ));
  assign new_n203_ = (~new_n205_ | (\a[5]  ^ (new_n204_ & (~new_n50_ | ~new_n201_)))) & ((~new_n206_ & (new_n207_ | ~new_n208_)) | (new_n205_ & (~\a[5]  ^ (new_n204_ & (~new_n50_ | ~new_n201_)))) | (~new_n205_ & (~\a[5]  | ~new_n204_ | (new_n50_ & new_n201_)) & (\a[5]  | (new_n204_ & (~new_n50_ | ~new_n201_)))));
  assign new_n204_ = (~\b[3]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[4]  | (~\a[4]  ^ ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[2]  | (~\a[3]  ^ ~\a[4] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  ^ ~\a[3] ));
  assign new_n205_ = ((\b[0]  & (\a[5]  ^ ~\a[6] ) & (\a[6]  | \a[7] ) & (~\a[6]  | ~\a[7] )) | (\b[1]  & (\a[7]  ^ ~\a[8] ) & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] )) | ((\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] ) & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (\b[0]  ^ \b[1] ))) ^ (\a[8]  & \b[0]  & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ));
  assign new_n206_ = \b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (~\b[0]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[4]  ^ ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\b[0]  ^ \b[1] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[4]  ^ ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[1]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  ^ ~\a[3] ));
  assign new_n207_ = \a[5]  ^ (((~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | (~\a[4]  ^ ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[2]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[3]  ^ ~\a[4] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n208_ = (\b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] )) ^ ((~\b[0]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[4]  ^ ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\b[0]  ^ \b[1] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[2]  | (~\a[4]  ^ ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[1]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n209_ = (~\a[8]  | ((~\b[0]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[7]  ^ ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\b[0]  ^ \b[1] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )))) ^ ((~\b[1]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[2]  | (~\a[7]  ^ ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n210_ = \a[5]  ^ (((\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\b[9]  ^ ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))))))) & (~\b[9]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[8]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n211_ = \a[5]  ^ (((\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n60_ & (~\b[7]  ^ \b[8] ))) & (~\b[7]  | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[8]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[6]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n212_ = ~new_n188_ ^ (~new_n126_ ^ new_n187_);
  assign new_n213_ = \a[5]  ^ ((new_n118_ ^ \a[8] ) ^ (new_n119_ | (~new_n121_ & new_n143_)));
  assign new_n214_ = \a[8]  ^ (~new_n215_ ^ new_n216_);
  assign new_n215_ = (~\a[11]  | (((new_n36_ & \a[14] ) | (~new_n70_ & (~new_n36_ | ~\a[14] ) & (new_n36_ | \a[14] ))) & (~\a[14]  | (~new_n153_ & new_n154_) | (new_n153_ & ~new_n154_)) & (\a[14]  | (~new_n153_ ^ new_n154_))) | ((~new_n36_ | ~\a[14] ) & (new_n70_ | (new_n36_ & \a[14] ) | (~new_n36_ & ~\a[14] )) & (~\a[14]  ^ (~new_n153_ ^ new_n154_)))) & (((~\a[11]  | (~new_n70_ & (~new_n36_ | ~\a[14] ) & (new_n36_ | \a[14] )) | (new_n70_ & (~new_n36_ ^ \a[14] ))) & (((~new_n157_ | ~\a[11] ) & (new_n163_ | (new_n157_ & \a[11] ) | (~new_n157_ & ~\a[11] ))) | (\a[11]  & (new_n70_ | (new_n36_ & \a[14] ) | (~new_n36_ & ~\a[14] )) & (~new_n70_ | (new_n36_ ^ \a[14] ))) | (~\a[11]  & (new_n70_ ^ (new_n36_ ^ \a[14] ))))) | (\a[11]  & (((~new_n36_ | ~\a[14] ) & (new_n70_ | (new_n36_ & \a[14] ) | (~new_n36_ & ~\a[14] ))) | (\a[14]  & (new_n153_ | ~new_n154_) & (~new_n153_ | new_n154_)) | (~\a[14]  & (new_n153_ ^ new_n154_))) & ((new_n36_ & \a[14] ) | (~new_n70_ & (~new_n36_ | ~\a[14] ) & (new_n36_ | \a[14] )) | (\a[14]  ^ (~new_n153_ ^ new_n154_)))) | (~\a[11]  & (((~new_n36_ | ~\a[14] ) & (new_n70_ | (new_n36_ & \a[14] ) | (~new_n36_ & ~\a[14] ))) ^ (\a[14]  ^ (~new_n153_ ^ new_n154_)))));
  assign new_n216_ = \a[11]  ^ (~new_n217_ ^ ((~\a[14]  | (new_n153_ & ~new_n154_) | (~new_n153_ & new_n154_)) & (((~new_n36_ | ~\a[14] ) & (new_n70_ | (new_n36_ & \a[14] ) | (~new_n36_ & ~\a[14] ))) | (\a[14]  & (~new_n153_ | new_n154_) & (new_n153_ | ~new_n154_)) | (~\a[14]  & (~new_n153_ ^ ~new_n154_)))));
  assign new_n217_ = \a[14]  ^ (~new_n218_ ^ new_n219_);
  assign new_n218_ = (new_n155_ | new_n156_) & ((new_n155_ & new_n156_) | (~new_n155_ & ~new_n156_) | ((new_n65_ | new_n67_) & (((new_n68_ | new_n69_) & ((new_n68_ & new_n69_) | (~new_n68_ & ~new_n69_) | (~new_n38_ & ~new_n63_))) | (~new_n65_ & ~new_n67_) | (new_n65_ & new_n67_))));
  assign new_n219_ = \a[17]  ? ((~\a[18]  | ~\b[8] ) & (~\b[9]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] ))) : (\a[18]  & \b[9] );
  assign new_n220_ = (~\a[8]  | ((~new_n152_ | ~\a[11] ) & (new_n152_ | \a[11] ) & ((new_n35_ & \a[11] ) | (((new_n157_ & \a[11] ) | (((new_n158_ & \a[11] ) | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] ))) & (~new_n157_ | ~\a[11] ) & (new_n157_ | \a[11] ))) & (~new_n35_ | ~\a[11] ) & (new_n35_ | \a[11] )))) | ((~new_n152_ ^ \a[11] ) & (~new_n35_ | ~\a[11] ) & (((~new_n157_ | ~\a[11] ) & (((~new_n158_ | ~\a[11] ) & (new_n160_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] ))) | (new_n157_ & \a[11] ) | (~new_n157_ & ~\a[11] ))) | (new_n35_ & \a[11] ) | (~new_n35_ & ~\a[11] )))) & (((~\a[8]  | (((new_n157_ & \a[11] ) | (((new_n158_ & \a[11] ) | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] ))) & (~new_n157_ | ~\a[11] ) & (new_n157_ | \a[11] ))) & (~new_n35_ | ~\a[11] ) & (new_n35_ | \a[11] )) | ((~new_n157_ | ~\a[11] ) & (((~new_n158_ | ~\a[11] ) & (new_n160_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] ))) | (new_n157_ & \a[11] ) | (~new_n157_ & ~\a[11] )) & (~new_n35_ ^ \a[11] ))) & (((~\a[8]  | (((new_n158_ & \a[11] ) | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] ))) & (~new_n157_ | ~\a[11] ) & (new_n157_ | \a[11] )) | ((~new_n158_ | ~\a[11] ) & (new_n160_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] )) & (~new_n157_ ^ \a[11] ))) & (((~\a[8]  | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] )) | (new_n160_ & (~new_n158_ ^ \a[11] ))) & (new_n95_ | (\a[8]  & (new_n160_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] )) & (~new_n160_ | (new_n158_ ^ \a[11] ))) | (~\a[8]  & (new_n160_ ^ (new_n158_ ^ \a[11] ))))) | (\a[8]  & (((~new_n158_ | ~\a[11] ) & (new_n160_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] ))) | (new_n157_ & \a[11] ) | (~new_n157_ & ~\a[11] )) & ((new_n158_ & \a[11] ) | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] )) | (new_n157_ ^ \a[11] ))) | (~\a[8]  & (((~new_n158_ | ~\a[11] ) & (new_n160_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] ))) ^ (new_n157_ ^ \a[11] ))))) | (\a[8]  & (((~new_n157_ | ~\a[11] ) & (((~new_n158_ | ~\a[11] ) & (new_n160_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] ))) | (new_n157_ & \a[11] ) | (~new_n157_ & ~\a[11] ))) | (new_n35_ & \a[11] ) | (~new_n35_ & ~\a[11] )) & ((new_n157_ & \a[11] ) | (((new_n158_ & \a[11] ) | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] ))) & (~new_n157_ | ~\a[11] ) & (new_n157_ | \a[11] )) | (new_n35_ ^ \a[11] ))) | (~\a[8]  & (((~new_n157_ | ~\a[11] ) & (((~new_n158_ | ~\a[11] ) & (new_n160_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] ))) | (new_n157_ & \a[11] ) | (~new_n157_ & ~\a[11] ))) ^ (new_n35_ ^ \a[11] ))))) | (\a[8]  & ((new_n152_ & \a[11] ) | (~new_n152_ & ~\a[11] ) | ((~new_n35_ | ~\a[11] ) & (((~new_n157_ | ~\a[11] ) & (((~new_n158_ | ~\a[11] ) & (new_n160_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] ))) | (new_n157_ & \a[11] ) | (~new_n157_ & ~\a[11] ))) | (new_n35_ & \a[11] ) | (~new_n35_ & ~\a[11] )))) & ((new_n152_ ^ \a[11] ) | (new_n35_ & \a[11] ) | (((new_n157_ & \a[11] ) | (((new_n158_ & \a[11] ) | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] ))) & (~new_n157_ | ~\a[11] ) & (new_n157_ | \a[11] ))) & (~new_n35_ | ~\a[11] ) & (new_n35_ | \a[11] )))) | (~\a[8]  & ((~new_n152_ ^ \a[11] ) ^ ((new_n35_ & \a[11] ) | (((new_n157_ & \a[11] ) | (((new_n158_ & \a[11] ) | (~new_n160_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] ))) & (~new_n157_ | ~\a[11] ) & (new_n157_ | \a[11] ))) & (~new_n35_ | ~\a[11] ) & (new_n35_ | \a[11] ))))));
  assign new_n221_ = (~\a[2]  | ((~new_n34_ | ~\a[5] ) & (new_n34_ | \a[5] ) & ((new_n161_ & \a[5] ) | (~new_n171_ & (new_n161_ | \a[5] ) & (~new_n161_ | ~\a[5] )))) | ((~new_n34_ ^ \a[5] ) & (~new_n161_ | ~\a[5] ) & (new_n171_ | (~new_n161_ & ~\a[5] ) | (new_n161_ & \a[5] )))) & (((~\a[2]  | (~new_n171_ & (new_n161_ | \a[5] ) & (~new_n161_ | ~\a[5] )) | (new_n171_ & (new_n161_ ^ ~\a[5] ))) & (((~new_n222_ | ~\a[2] ) & (new_n223_ | (new_n222_ & \a[2] ) | (~new_n222_ & ~\a[2] ))) | (\a[2]  & (new_n171_ | (~new_n161_ & ~\a[5] ) | (new_n161_ & \a[5] )) & (~new_n171_ | (~new_n161_ ^ ~\a[5] ))) | (~\a[2]  & (new_n171_ ^ (~new_n161_ ^ ~\a[5] ))))) | (\a[2]  & ((new_n34_ & \a[5] ) | (~new_n34_ & ~\a[5] ) | ((~new_n161_ | ~\a[5] ) & (new_n171_ | (~new_n161_ & ~\a[5] ) | (new_n161_ & \a[5] )))) & ((new_n34_ ^ \a[5] ) | (new_n161_ & \a[5] ) | (~new_n171_ & (new_n161_ | \a[5] ) & (~new_n161_ | ~\a[5] )))) | (~\a[2]  & ((~new_n34_ ^ \a[5] ) ^ ((new_n161_ & \a[5] ) | (~new_n171_ & (new_n161_ | \a[5] ) & (~new_n161_ | ~\a[5] ))))));
  assign new_n222_ = ((new_n172_ & \a[5] ) | (((new_n173_ & \a[5] ) | (~new_n174_ & (~new_n173_ | ~\a[5] ) & (new_n173_ | \a[5] ))) & (~new_n172_ | ~\a[5] ) & (new_n172_ | \a[5] ))) ^ (\a[5]  ^ (~new_n165_ ^ new_n169_));
  assign new_n223_ = (~\a[2]  | ((~new_n172_ | ~\a[5] ) & (new_n172_ | \a[5] ) & ((new_n173_ & \a[5] ) | ((~new_n173_ | ~\a[5] ) & (new_n173_ | \a[5] ) & ((new_n224_ & \a[5] ) | ((~new_n224_ | ~\a[5] ) & (new_n224_ | \a[5] ) & ((new_n178_ & \a[5] ) | (~new_n225_ & (~new_n178_ | ~\a[5] ) & (new_n178_ | \a[5] )))))))) | ((~new_n172_ ^ \a[5] ) & (~new_n173_ | ~\a[5] ) & ((new_n173_ & \a[5] ) | (~new_n173_ & ~\a[5] ) | ((~new_n224_ | ~\a[5] ) & ((new_n224_ & \a[5] ) | (~new_n224_ & ~\a[5] ) | ((~new_n178_ | ~\a[5] ) & (new_n225_ | (new_n178_ & \a[5] ) | (~new_n178_ & ~\a[5] )))))))) & (((~\a[2]  | ((~new_n173_ | ~\a[5] ) & (new_n173_ | \a[5] ) & ((new_n224_ & \a[5] ) | ((~new_n224_ | ~\a[5] ) & (new_n224_ | \a[5] ) & ((new_n178_ & \a[5] ) | (~new_n225_ & (~new_n178_ | ~\a[5] ) & (new_n178_ | \a[5] )))))) | ((~new_n173_ ^ \a[5] ) & (~new_n224_ | ~\a[5] ) & ((new_n224_ & \a[5] ) | (~new_n224_ & ~\a[5] ) | ((~new_n178_ | ~\a[5] ) & (new_n225_ | (new_n178_ & \a[5] ) | (~new_n178_ & ~\a[5] )))))) & (((~\a[2]  | ((~new_n224_ | ~\a[5] ) & (new_n224_ | \a[5] ) & ((new_n178_ & \a[5] ) | (~new_n225_ & (~new_n178_ | ~\a[5] ) & (new_n178_ | \a[5] )))) | ((~new_n224_ ^ \a[5] ) & (~new_n178_ | ~\a[5] ) & (new_n225_ | (new_n178_ & \a[5] ) | (~new_n178_ & ~\a[5] )))) & (((~\a[2]  | (~new_n225_ & (~new_n178_ | ~\a[5] ) & (new_n178_ | \a[5] )) | (new_n225_ & (~new_n178_ ^ \a[5] ))) & (new_n227_ | (\a[2]  & (new_n225_ | (new_n178_ & \a[5] ) | (~new_n178_ & ~\a[5] )) & (~new_n225_ | (new_n178_ ^ \a[5] ))) | (~\a[2]  & (new_n225_ ^ (new_n178_ ^ \a[5] ))))) | (\a[2]  & ((new_n224_ & \a[5] ) | (~new_n224_ & ~\a[5] ) | ((~new_n178_ | ~\a[5] ) & (new_n225_ | (new_n178_ & \a[5] ) | (~new_n178_ & ~\a[5] )))) & ((new_n224_ ^ \a[5] ) | (new_n178_ & \a[5] ) | (~new_n225_ & (~new_n178_ | ~\a[5] ) & (new_n178_ | \a[5] )))) | (~\a[2]  & ((~new_n224_ ^ \a[5] ) ^ ((new_n178_ & \a[5] ) | (~new_n225_ & (~new_n178_ | ~\a[5] ) & (new_n178_ | \a[5] ))))))) | (\a[2]  & ((new_n173_ & \a[5] ) | (~new_n173_ & ~\a[5] ) | ((~new_n224_ | ~\a[5] ) & ((new_n224_ & \a[5] ) | (~new_n224_ & ~\a[5] ) | ((~new_n178_ | ~\a[5] ) & (new_n225_ | (new_n178_ & \a[5] ) | (~new_n178_ & ~\a[5] )))))) & ((new_n173_ ^ \a[5] ) | (new_n224_ & \a[5] ) | ((~new_n224_ | ~\a[5] ) & (new_n224_ | \a[5] ) & ((new_n178_ & \a[5] ) | (~new_n225_ & (~new_n178_ | ~\a[5] ) & (new_n178_ | \a[5] )))))) | (~\a[2]  & ((~new_n173_ ^ \a[5] ) ^ ((new_n224_ & \a[5] ) | ((~new_n224_ | ~\a[5] ) & (new_n224_ | \a[5] ) & ((new_n178_ & \a[5] ) | (~new_n225_ & (~new_n178_ | ~\a[5] ) & (new_n178_ | \a[5] ))))))))) | (\a[2]  & ((new_n172_ & \a[5] ) | (~new_n172_ & ~\a[5] ) | ((~new_n173_ | ~\a[5] ) & ((new_n173_ & \a[5] ) | (~new_n173_ & ~\a[5] ) | ((~new_n224_ | ~\a[5] ) & ((new_n224_ & \a[5] ) | (~new_n224_ & ~\a[5] ) | ((~new_n178_ | ~\a[5] ) & (new_n225_ | (new_n178_ & \a[5] ) | (~new_n178_ & ~\a[5] )))))))) & ((new_n172_ ^ \a[5] ) | (new_n173_ & \a[5] ) | ((~new_n173_ | ~\a[5] ) & (new_n173_ | \a[5] ) & ((new_n224_ & \a[5] ) | ((~new_n224_ | ~\a[5] ) & (new_n224_ | \a[5] ) & ((new_n178_ & \a[5] ) | (~new_n225_ & (~new_n178_ | ~\a[5] ) & (new_n178_ | \a[5] )))))))) | (~\a[2]  & ((~new_n172_ ^ \a[5] ) ^ ((new_n173_ & \a[5] ) | ((~new_n173_ | ~\a[5] ) & (new_n173_ | \a[5] ) & ((new_n224_ & \a[5] ) | ((~new_n224_ | ~\a[5] ) & (new_n224_ | \a[5] ) & ((new_n178_ & \a[5] ) | (~new_n225_ & (~new_n178_ | ~\a[5] ) & (new_n178_ | \a[5] ))))))))));
  assign new_n224_ = ~new_n175_ ^ new_n177_;
  assign new_n225_ = (~new_n179_ | ~\a[5] ) & (~new_n226_ | (~new_n180_ & (new_n181_ | ~new_n213_)));
  assign new_n226_ = \a[5]  ^ ((new_n97_ ^ \a[8] ) ^ ((new_n118_ & \a[8] ) | ((new_n119_ | (~new_n121_ & new_n143_)) & (new_n118_ | \a[8] ) & (~new_n118_ | ~\a[8] ))));
  assign new_n227_ = (~\a[2]  | (new_n226_ & (new_n180_ | (~new_n181_ & new_n213_))) | (~new_n226_ & ~new_n180_ & (new_n181_ | ~new_n213_))) & (((~\a[2]  | (~new_n181_ & new_n213_) | (new_n181_ & ~new_n213_)) & (((~new_n228_ | ~\a[2] ) & ((new_n228_ & \a[2] ) | (~new_n228_ & ~\a[2] ) | ((~new_n229_ | ~\a[2] ) & (new_n230_ | (new_n229_ & \a[2] ) | (~new_n229_ & ~\a[2] ))))) | (\a[2]  & (new_n181_ | ~new_n213_) & (~new_n181_ | new_n213_)) | (~\a[2]  & (new_n181_ ^ new_n213_)))) | (\a[2]  & (~new_n226_ | (~new_n180_ & (new_n181_ | ~new_n213_))) & (new_n226_ | new_n180_ | (~new_n181_ & new_n213_))) | (~\a[2]  & (~new_n226_ ^ (new_n180_ | (~new_n181_ & new_n213_)))));
  assign new_n228_ = (\a[5]  ^ (~new_n121_ ^ new_n143_)) ^ ((new_n182_ & \a[5] ) | ((~new_n182_ | ~\a[5] ) & (new_n182_ | \a[5] ) & ((new_n185_ & \a[5] ) | ((~new_n185_ | ~\a[5] ) & (new_n185_ | \a[5] ) & (new_n186_ | (~new_n189_ & new_n212_))))));
  assign new_n229_ = (new_n182_ ^ \a[5] ) ^ ((new_n185_ & \a[5] ) | ((new_n185_ | \a[5] ) & (~new_n185_ | ~\a[5] ) & ((~new_n188_ & (new_n126_ | ~new_n187_) & (~new_n126_ | new_n187_)) | (~new_n189_ & (new_n188_ | (~new_n126_ & new_n187_) | (new_n126_ & ~new_n187_)) & (~new_n188_ | (~new_n126_ ^ new_n187_))))));
  assign new_n230_ = (~\a[2]  | (new_n231_ & (new_n186_ | (~new_n189_ & new_n212_))) | (~new_n231_ & ~new_n186_ & (new_n189_ | ~new_n212_))) & (((~\a[2]  | (~new_n189_ & new_n212_) | (new_n189_ & ~new_n212_)) & (((~new_n232_ | ~\a[2] ) & ((new_n232_ & \a[2] ) | (~new_n232_ & ~\a[2] ) | ((~new_n234_ | ~\a[2] ) & (new_n235_ | (new_n234_ & \a[2] ) | (~new_n234_ & ~\a[2] ))))) | (\a[2]  & (new_n189_ | ~new_n212_) & (~new_n189_ | new_n212_)) | (~\a[2]  & (new_n189_ ^ new_n212_)))) | (\a[2]  & (~new_n231_ | (~new_n186_ & (new_n189_ | ~new_n212_))) & (new_n231_ | new_n186_ | (~new_n189_ & new_n212_))) | (~\a[2]  & (~new_n231_ ^ (new_n186_ | (~new_n189_ & new_n212_)))));
  assign new_n231_ = \a[5]  ^ (((~new_n142_ & (new_n106_ | (~new_n105_ & new_n113_) | (new_n105_ & ~new_n113_)) & (~new_n106_ | (~new_n105_ ^ new_n113_))) | (~new_n126_ & (new_n142_ | (~new_n106_ & (new_n105_ | ~new_n113_) & (~new_n105_ | new_n113_)) | (new_n106_ & (new_n105_ ^ new_n113_))) & (~new_n142_ | (~new_n106_ ^ (~new_n105_ ^ new_n113_))))) ^ (~new_n125_ ^ (new_n183_ ^ ((~new_n105_ & new_n113_) | (~new_n106_ & (new_n105_ | ~new_n113_) & (~new_n105_ | new_n113_))))));
  assign new_n232_ = new_n233_ ^ (new_n192_ | (~new_n192_ & ~new_n194_ & ((~new_n211_ & (new_n132_ | (~new_n131_ & new_n139_) | (new_n131_ & ~new_n139_)) & (~new_n132_ | (~new_n131_ ^ new_n139_))) | (~new_n195_ & (new_n211_ | (~new_n132_ & (new_n131_ | ~new_n139_) & (~new_n131_ | new_n139_)) | (new_n132_ & (new_n131_ ^ new_n139_))) & (~new_n211_ | (~new_n132_ ^ (~new_n131_ ^ new_n139_)))))));
  assign new_n233_ = ~new_n210_ ^ ((~new_n127_ ^ new_n128_) ^ ((new_n129_ & ~new_n130_) | ((new_n129_ | ~new_n130_) & (~new_n129_ | new_n130_) & ((~new_n131_ & new_n139_) | (~new_n132_ & (new_n131_ | ~new_n139_) & (~new_n131_ | new_n139_))))));
  assign new_n234_ = (~new_n192_ & ~new_n194_) ^ ((~new_n211_ & (new_n132_ | (~new_n131_ & new_n139_) | (new_n131_ & ~new_n139_)) & (~new_n132_ | (~new_n131_ ^ new_n139_))) | (~new_n195_ & (new_n211_ | (~new_n132_ & (new_n131_ | ~new_n139_) & (~new_n131_ | new_n139_)) | (new_n132_ & (new_n131_ ^ new_n139_))) & (~new_n211_ | (~new_n132_ ^ (~new_n131_ ^ new_n139_)))));
  assign new_n235_ = (new_n237_ | (~new_n195_ & new_n236_) | (new_n195_ & ~new_n236_)) & ((~new_n237_ & (new_n195_ | ~new_n236_) & (~new_n195_ | new_n236_)) | (new_n237_ & (new_n195_ ^ new_n236_)) | ((~new_n238_ | new_n256_) & ((~new_n239_ & (new_n241_ | ~new_n255_)) | (~new_n238_ & new_n256_) | (new_n238_ & ~new_n256_))));
  assign new_n236_ = ~new_n211_ ^ (~new_n132_ ^ (~new_n131_ ^ new_n139_));
  assign new_n237_ = \a[2]  ^ (~\b[9]  | ((new_n66_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & ((~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] )));
  assign new_n238_ = (~new_n196_ ^ new_n197_) ^ ((new_n198_ & ~new_n199_) | ((new_n198_ | ~new_n199_) & (~new_n198_ | new_n199_) & ((~new_n200_ & new_n209_) | (~new_n203_ & (new_n200_ | ~new_n209_) & (~new_n200_ | new_n209_)))));
  assign new_n239_ = ~new_n240_ & ((~new_n198_ & new_n199_) | (new_n198_ & ~new_n199_) | ((new_n200_ | ~new_n209_) & (new_n203_ | (~new_n200_ & new_n209_) | (new_n200_ & ~new_n209_)))) & ((~new_n198_ ^ new_n199_) | (~new_n200_ & new_n209_) | (~new_n203_ & (new_n200_ | ~new_n209_) & (~new_n200_ | new_n209_)));
  assign new_n240_ = \a[2]  ^ ((~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )))) | ((~\b[8]  ^ \b[9] ) & (~\b[7]  | ~\b[8] ) & (new_n60_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )))) & (~\b[7]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[9]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[8]  | \a[0]  | ~\a[1] ));
  assign new_n241_ = (new_n243_ | (~new_n203_ & new_n242_) | (new_n203_ & ~new_n242_)) & ((~new_n243_ & (new_n203_ | ~new_n242_) & (~new_n203_ | new_n242_)) | (new_n243_ & (new_n203_ ^ new_n242_)) | ((new_n244_ | ~new_n245_) & ((~new_n244_ & new_n245_) | (new_n244_ & ~new_n245_) | ((new_n246_ | ~new_n247_) & (new_n248_ | (~new_n246_ & new_n247_) | (new_n246_ & ~new_n247_))))));
  assign new_n242_ = new_n209_ ^ (~\a[5]  ^ (new_n202_ & (~new_n47_ | ~new_n201_)));
  assign new_n243_ = \a[2]  ^ ((~\b[6]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[8]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[7]  | \a[0]  | ~\a[1] ) & ((~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n60_ & (~\b[7]  ^ \b[8] )) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )));
  assign new_n244_ = \a[2]  ^ ((~\b[5]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[7]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[6]  | \a[0]  | ~\a[1] ) & (~new_n41_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )));
  assign new_n245_ = (new_n206_ | (~new_n207_ & new_n208_)) ^ (new_n205_ ^ (~\a[5]  ^ (new_n204_ & (~new_n50_ | ~new_n201_))));
  assign new_n246_ = \a[2]  ^ ((~\b[4]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[6]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[5]  | \a[0]  | ~\a[1] ) & (~new_n44_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )));
  assign new_n247_ = ~new_n207_ ^ new_n208_;
  assign new_n248_ = (~new_n251_ | (\a[2]  ^ (new_n250_ & (~new_n47_ | ~new_n249_)))) & ((new_n251_ & (~\a[2]  ^ (new_n250_ & (~new_n47_ | ~new_n249_)))) | (~new_n251_ & (~\a[2]  | ~new_n250_ | (new_n47_ & new_n249_)) & (\a[2]  | (new_n250_ & (~new_n47_ | ~new_n249_)))) | ((new_n252_ | ~new_n253_) & (new_n254_ | (~new_n252_ & new_n253_) | (new_n252_ & ~new_n253_))));
  assign new_n249_ = \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] );
  assign new_n250_ = (~\b[3]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[5]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[4]  | \a[0]  | ~\a[1] );
  assign new_n251_ = (~\a[5]  | ((~\b[0]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[4]  ^ ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\b[0]  ^ \b[1] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )))) ^ ((~\b[1]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[2]  | (~\a[4]  ^ ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\b[2]  ^ (\b[0]  | ~\b[1] ))) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n252_ = \a[2]  ^ ((~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )))) | ((~\b[3]  ^ \b[4] ) & (~\b[2]  | ~\b[3] ) & ((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[4]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[3]  | \a[0]  | ~\a[1] ));
  assign new_n253_ = ((\b[0]  & (\a[2]  ^ ~\a[3] ) & (\a[3]  | \a[4] ) & (~\a[3]  | ~\a[4] )) | (\b[1]  & (\a[4]  ^ ~\a[5] ) & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] )) | ((\a[4]  | \a[5] ) & (~\a[4]  | ~\a[5] ) & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (\b[0]  ^ \b[1] ))) ^ (\a[5]  & \b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ));
  assign new_n254_ = (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[2]  ^ ((((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] )))) & ((\b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (~\a[2]  ^ ((((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] )))) | ((~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\a[2]  | (((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )) & ((\b[2]  ^ \b[3] ) | (\b[1]  & (\b[0]  | \b[2] ))) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[3]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[1]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[2]  & ~\a[0]  & \a[1] )) & (\a[2]  | ((((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] )))) | (\b[2]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[1]  & ~\a[0]  & \a[1] ) | (\b[0]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | ((~\b[2]  ^ (\b[0]  | ~\b[1] )) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[0]  & ~\a[0]  & \a[1] ) | (\b[1]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | ((\b[0]  ^ \b[1] ) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | ~\a[2]  | (\a[0]  & \b[0] ));
  assign new_n255_ = ~new_n240_ ^ ((~new_n198_ ^ new_n199_) ^ ((~new_n200_ & new_n209_) | (~new_n203_ & (new_n200_ | ~new_n209_) & (~new_n200_ | new_n209_))));
  assign new_n256_ = \a[2]  ^ ((~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | (~\b[9]  ^ ((\b[8]  & \b[9] ) | ((~\b[8]  | ~\b[9] ) & (\b[8]  | \b[9] ) & ((\b[7]  & \b[8] ) | (~new_n60_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))))))) & (~\b[8]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | \a[0]  | \a[1] ) & (~\b[9]  | \a[0]  | ~\a[1] ));
  assign new_n257_ = new_n258_ ^ (((~\a[5]  | (~new_n214_ & new_n220_) | (new_n214_ & ~new_n220_)) & (((~new_n34_ | ~\a[5] ) & ((new_n34_ & \a[5] ) | (~new_n34_ & ~\a[5] ) | ((~new_n161_ | ~\a[5] ) & (new_n171_ | (~new_n161_ & ~\a[5] ) | (new_n161_ & \a[5] ))))) | (\a[5]  & (new_n214_ | ~new_n220_) & (~new_n214_ | new_n220_)) | (~\a[5]  & (new_n214_ ^ new_n220_)))) ^ (~\a[5]  ^ ~\a[14] ));
  assign new_n258_ = ((~new_n259_ | ~\a[11] ) & (new_n215_ | (~new_n259_ & ~\a[11] ) | (new_n259_ & \a[11] ))) ^ (~\a[17]  | (\a[18]  & \b[9] ));
  assign new_n259_ = ~new_n217_ ^ ((~\a[14]  | (new_n153_ & ~new_n154_) | (~new_n153_ & new_n154_)) & (((~new_n36_ | ~\a[14] ) & (new_n70_ | (new_n36_ & \a[14] ) | (~new_n36_ & ~\a[14] ))) | (\a[14]  & (~new_n153_ | new_n154_) & (new_n153_ | ~new_n154_)) | (~\a[14]  & (~new_n153_ ^ ~new_n154_))));
  assign new_n260_ = (new_n261_ ^ ((\a[8]  & (new_n215_ | ~new_n216_) & (~new_n215_ | new_n216_)) | (~new_n220_ & (~\a[8]  | (~new_n215_ & new_n216_) | (new_n215_ & ~new_n216_)) & (\a[8]  | (~new_n215_ ^ new_n216_))))) ^ (new_n262_ ^ (\a[2]  ^ \a[8] ));
  assign new_n261_ = (~\a[14]  | (~new_n218_ & new_n219_) | (new_n218_ & ~new_n219_)) & (((~\a[14]  | (~new_n153_ & new_n154_) | (new_n153_ & ~new_n154_)) & (((~new_n36_ | ~\a[14] ) & (new_n70_ | (new_n36_ & \a[14] ) | (~new_n36_ & ~\a[14] ))) | (\a[14]  & (new_n153_ | ~new_n154_) & (~new_n153_ | new_n154_)) | (~\a[14]  & (new_n153_ ^ new_n154_)))) | (\a[14]  & (new_n218_ | ~new_n219_) & (~new_n218_ | new_n219_)) | (~\a[14]  & (new_n218_ ^ new_n219_)));
  assign new_n262_ = \a[11]  ^ ((\a[17]  & ((\a[18]  & \b[8] ) | (\b[9]  & (\a[17]  | \a[18] ) & (~\a[17]  | ~\a[18] )))) | (~new_n218_ & (~\a[17]  | ((~\a[18]  | ~\b[8] ) & (~\b[9]  | (~\a[17]  & ~\a[18] ) | (\a[17]  & \a[18] )))) & (\a[17]  | (\a[18]  & \b[9] ))));
  assign new_n263_ = ((\a[2]  & (new_n171_ | (~new_n161_ & ~\a[5] ) | (new_n161_ & \a[5] )) & (~new_n171_ | (~new_n161_ ^ ~\a[5] ))) | (((new_n222_ & \a[2] ) | (~new_n223_ & (~new_n222_ | ~\a[2] ) & (new_n222_ | \a[2] ))) & (~\a[2]  | (~new_n171_ & (new_n161_ | \a[5] ) & (~new_n161_ | ~\a[5] )) | (new_n171_ & (new_n161_ ^ ~\a[5] ))) & (\a[2]  | (~new_n171_ ^ (~new_n161_ ^ ~\a[5] ))))) ^ (\a[2]  ^ ((new_n34_ ^ \a[5] ) ^ ((new_n161_ & \a[5] ) | (~new_n171_ & (new_n161_ | \a[5] ) & (~new_n161_ | ~\a[5] )))));
  assign new_n264_ = ((~new_n265_ ^ \a[2] ) ^ ((new_n222_ & \a[2] ) | ((~new_n222_ | ~\a[2] ) & (new_n222_ | \a[2] ) & ((new_n266_ & \a[2] ) | (~new_n267_ & (~new_n266_ | ~\a[2] ) & (new_n266_ | \a[2] )))))) & ((~new_n222_ ^ \a[2] ) ^ ((new_n266_ & \a[2] ) | (~new_n267_ & (~new_n266_ | ~\a[2] ) & (new_n266_ | \a[2] )))) & (new_n267_ ^ (new_n266_ ^ \a[2] )) & ~new_n268_ & ~new_n269_ & new_n270_;
  assign new_n265_ = ((\a[5]  & (new_n165_ | ~new_n169_) & (~new_n165_ | new_n169_)) | (((new_n172_ & \a[5] ) | ((~new_n172_ | ~\a[5] ) & (new_n172_ | \a[5] ) & ((new_n173_ & \a[5] ) | (~new_n174_ & (~new_n173_ | ~\a[5] ) & (new_n173_ | \a[5] ))))) & (~\a[5]  | (~new_n165_ & new_n169_) | (new_n165_ & ~new_n169_)) & (\a[5]  | (~new_n165_ ^ new_n169_)))) ^ (\a[5]  ^ (new_n170_ ^ (new_n162_ | (~new_n165_ & new_n169_))));
  assign new_n266_ = ((new_n173_ & \a[5] ) | (~new_n174_ & (~new_n173_ | ~\a[5] ) & (new_n173_ | \a[5] ))) ^ (~new_n172_ ^ ~\a[5] );
  assign new_n267_ = (~\a[2]  | ((~new_n173_ | ~\a[5] ) & (new_n173_ | \a[5] ) & ((new_n224_ & \a[5] ) | ((new_n224_ | \a[5] ) & (~new_n224_ | ~\a[5] ) & ((new_n178_ & \a[5] ) | (~new_n225_ & (new_n178_ | \a[5] ) & (~new_n178_ | ~\a[5] )))))) | ((~new_n173_ ^ \a[5] ) & (~new_n224_ | ~\a[5] ) & ((~new_n224_ & ~\a[5] ) | (new_n224_ & \a[5] ) | ((~new_n178_ | ~\a[5] ) & (new_n225_ | (~new_n178_ & ~\a[5] ) | (new_n178_ & \a[5] )))))) & (((~\a[2]  | ((new_n224_ | \a[5] ) & (~new_n224_ | ~\a[5] ) & ((new_n178_ & \a[5] ) | (~new_n225_ & (new_n178_ | \a[5] ) & (~new_n178_ | ~\a[5] )))) | ((new_n224_ ^ ~\a[5] ) & (~new_n178_ | ~\a[5] ) & (new_n225_ | (~new_n178_ & ~\a[5] ) | (new_n178_ & \a[5] )))) & (((~\a[2]  | (~new_n225_ & (new_n178_ | \a[5] ) & (~new_n178_ | ~\a[5] )) | (new_n225_ & (new_n178_ ^ ~\a[5] ))) & (new_n227_ | (\a[2]  & (new_n225_ | (~new_n178_ & ~\a[5] ) | (new_n178_ & \a[5] )) & (~new_n225_ | (~new_n178_ ^ ~\a[5] ))) | (~\a[2]  & (new_n225_ ^ (~new_n178_ ^ ~\a[5] ))))) | (\a[2]  & ((~new_n224_ & ~\a[5] ) | (new_n224_ & \a[5] ) | ((~new_n178_ | ~\a[5] ) & (new_n225_ | (~new_n178_ & ~\a[5] ) | (new_n178_ & \a[5] )))) & ((~new_n224_ ^ ~\a[5] ) | (new_n178_ & \a[5] ) | (~new_n225_ & (new_n178_ | \a[5] ) & (~new_n178_ | ~\a[5] )))) | (~\a[2]  & ((new_n224_ ^ ~\a[5] ) ^ ((new_n178_ & \a[5] ) | (~new_n225_ & (new_n178_ | \a[5] ) & (~new_n178_ | ~\a[5] ))))))) | (\a[2]  & ((new_n173_ & \a[5] ) | (~new_n173_ & ~\a[5] ) | ((~new_n224_ | ~\a[5] ) & ((~new_n224_ & ~\a[5] ) | (new_n224_ & \a[5] ) | ((~new_n178_ | ~\a[5] ) & (new_n225_ | (~new_n178_ & ~\a[5] ) | (new_n178_ & \a[5] )))))) & ((new_n173_ ^ \a[5] ) | (new_n224_ & \a[5] ) | ((new_n224_ | \a[5] ) & (~new_n224_ | ~\a[5] ) & ((new_n178_ & \a[5] ) | (~new_n225_ & (new_n178_ | \a[5] ) & (~new_n178_ | ~\a[5] )))))) | (~\a[2]  & ((~new_n173_ ^ \a[5] ) ^ ((new_n224_ & \a[5] ) | ((new_n224_ | \a[5] ) & (~new_n224_ | ~\a[5] ) & ((new_n178_ & \a[5] ) | (~new_n225_ & (new_n178_ | \a[5] ) & (~new_n178_ | ~\a[5] ))))))));
  assign new_n268_ = ((\a[2]  & ((~new_n224_ & ~\a[5] ) | (new_n224_ & \a[5] ) | ((~new_n178_ | ~\a[5] ) & (new_n225_ | (~new_n178_ & ~\a[5] ) | (new_n178_ & \a[5] )))) & ((~new_n224_ ^ ~\a[5] ) | (new_n178_ & \a[5] ) | (~new_n225_ & (new_n178_ | \a[5] ) & (~new_n178_ | ~\a[5] )))) | (((\a[2]  & (new_n225_ | (~new_n178_ & ~\a[5] ) | (new_n178_ & \a[5] )) & (~new_n225_ | (~new_n178_ ^ ~\a[5] ))) | (~new_n227_ & (~\a[2]  | (~new_n225_ & (new_n178_ | \a[5] ) & (~new_n178_ | ~\a[5] )) | (new_n225_ & (new_n178_ ^ ~\a[5] ))) & (\a[2]  | (~new_n225_ ^ (~new_n178_ ^ ~\a[5] ))))) & (~\a[2]  | ((new_n224_ | \a[5] ) & (~new_n224_ | ~\a[5] ) & ((new_n178_ & \a[5] ) | (~new_n225_ & (new_n178_ | \a[5] ) & (~new_n178_ | ~\a[5] )))) | ((new_n224_ ^ ~\a[5] ) & (~new_n178_ | ~\a[5] ) & (new_n225_ | (~new_n178_ & ~\a[5] ) | (new_n178_ & \a[5] )))) & (\a[2]  | ((~new_n224_ ^ ~\a[5] ) ^ ((new_n178_ & \a[5] ) | (~new_n225_ & (new_n178_ | \a[5] ) & (~new_n178_ | ~\a[5] ))))))) ^ (\a[2]  ^ ((new_n173_ ^ \a[5] ) ^ ((new_n224_ & \a[5] ) | ((new_n224_ | \a[5] ) & (~new_n224_ | ~\a[5] ) & ((new_n178_ & \a[5] ) | (~new_n225_ & (new_n178_ | \a[5] ) & (~new_n178_ | ~\a[5] )))))));
  assign new_n269_ = ((\a[2]  & (new_n225_ | (new_n178_ & \a[5] ) | (~new_n178_ & ~\a[5] )) & (~new_n225_ | (new_n178_ ^ \a[5] ))) | (~new_n227_ & (~\a[2]  | (~new_n225_ & (~new_n178_ | ~\a[5] ) & (new_n178_ | \a[5] )) | (new_n225_ & (~new_n178_ ^ \a[5] ))) & (\a[2]  | (~new_n225_ ^ (new_n178_ ^ \a[5] ))))) ^ (\a[2]  ^ ((new_n224_ ^ \a[5] ) ^ ((new_n178_ & \a[5] ) | (~new_n225_ & (~new_n178_ | ~\a[5] ) & (new_n178_ | \a[5] )))));
  assign new_n270_ = (((~new_n272_ | ~\a[2] ) & (new_n273_ | (new_n272_ & \a[2] ) | (~new_n272_ & ~\a[2] ))) ^ (\a[2]  ^ (~new_n225_ ^ new_n271_))) & (~new_n273_ | (new_n272_ ^ \a[2] )) & ~new_n274_ & new_n275_ & (new_n273_ | (new_n272_ & \a[2] ) | (~new_n272_ & ~\a[2] ));
  assign new_n271_ = ~new_n178_ ^ ~\a[5] ;
  assign new_n272_ = new_n226_ ^ (new_n180_ | (~new_n181_ & new_n213_));
  assign new_n273_ = (~\a[2]  | (~new_n181_ & new_n213_) | (new_n181_ & ~new_n213_)) & (((~new_n228_ | ~\a[2] ) & (((~new_n229_ | ~\a[2] ) & (new_n230_ | (new_n229_ & \a[2] ) | (~new_n229_ & ~\a[2] ))) | (new_n228_ & \a[2] ) | (~new_n228_ & ~\a[2] ))) | (\a[2]  & (new_n181_ | ~new_n213_) & (~new_n181_ | new_n213_)) | (~\a[2]  & (new_n181_ ^ new_n213_)));
  assign new_n274_ = ((new_n228_ & \a[2] ) | (((new_n229_ & \a[2] ) | (~new_n230_ & (~new_n229_ | ~\a[2] ) & (new_n229_ | \a[2] ))) & (~new_n228_ | ~\a[2] ) & (new_n228_ | \a[2] ))) ^ (\a[2]  ^ (~new_n181_ ^ new_n213_));
  assign new_n275_ = ((new_n228_ ^ \a[2] ) | (new_n229_ & \a[2] ) | (~new_n230_ & (~new_n229_ | ~\a[2] ) & (new_n229_ | \a[2] ))) & ((new_n228_ & \a[2] ) | (~new_n228_ & ~\a[2] ) | ((~new_n229_ | ~\a[2] ) & (new_n230_ | (new_n229_ & \a[2] ) | (~new_n229_ & ~\a[2] )))) & (new_n230_ ^ (new_n229_ ^ \a[2] )) & ~new_n277_ & ~new_n278_ & ~new_n276_ & new_n279_;
  assign new_n276_ = ((new_n232_ & \a[2] ) | (((new_n234_ & \a[2] ) | (~new_n235_ & (~new_n234_ | ~\a[2] ) & (new_n234_ | \a[2] ))) & (~new_n232_ | ~\a[2] ) & (new_n232_ | \a[2] ))) & (~\a[2]  | (~new_n189_ & new_n212_) | (new_n189_ & ~new_n212_)) & (\a[2]  | (~new_n189_ ^ new_n212_));
  assign new_n277_ = ((\a[2]  & (new_n189_ | ~new_n212_) & (~new_n189_ | new_n212_)) | (((new_n232_ & \a[2] ) | ((~new_n232_ | ~\a[2] ) & (new_n232_ | \a[2] ) & ((new_n234_ & \a[2] ) | (~new_n235_ & (~new_n234_ | ~\a[2] ) & (new_n234_ | \a[2] ))))) & (~\a[2]  | (~new_n189_ & new_n212_) | (new_n189_ & ~new_n212_)) & (\a[2]  | (~new_n189_ ^ new_n212_)))) ^ (\a[2]  ^ (new_n231_ ^ (new_n186_ | (~new_n189_ & new_n212_))));
  assign new_n278_ = (~new_n232_ | ~\a[2] ) & (((~new_n234_ | ~\a[2] ) & (new_n235_ | (new_n234_ & \a[2] ) | (~new_n234_ & ~\a[2] ))) | (new_n232_ & \a[2] ) | (~new_n232_ & ~\a[2] )) & (~\a[2]  ^ (~new_n189_ ^ new_n212_));
  assign new_n279_ = ((~new_n232_ ^ \a[2] ) ^ ((new_n234_ & \a[2] ) | (~new_n235_ & (new_n234_ | \a[2] ) & (~new_n234_ | ~\a[2] )))) & (new_n235_ ^ (~new_n234_ ^ ~\a[2] )) & (~new_n280_ | new_n281_) & new_n282_ & (new_n280_ | ~new_n281_);
  assign new_n280_ = (~new_n238_ | new_n256_) & ((~new_n239_ & (new_n241_ | ~new_n255_)) | (new_n238_ & ~new_n256_) | (~new_n238_ & new_n256_));
  assign new_n281_ = ~new_n237_ ^ (~new_n195_ ^ new_n236_);
  assign new_n282_ = (new_n285_ | new_n239_ | (~new_n241_ & new_n255_)) & (~new_n285_ | (~new_n239_ & (new_n241_ | ~new_n255_))) & (~new_n241_ | new_n255_) & (new_n241_ | ~new_n255_) & (~new_n283_ | new_n284_) & new_n286_ & (new_n283_ | ~new_n284_);
  assign new_n283_ = (new_n244_ | ~new_n245_) & ((~new_n244_ & new_n245_) | (new_n244_ & ~new_n245_) | ((new_n246_ | ~new_n247_) & (new_n248_ | (~new_n246_ & new_n247_) | (new_n246_ & ~new_n247_))));
  assign new_n284_ = ~new_n243_ ^ (~new_n203_ ^ new_n242_);
  assign new_n285_ = ~new_n256_ ^ ((~new_n196_ ^ new_n197_) ^ ((new_n198_ & ~new_n199_) | ((new_n198_ | ~new_n199_) & (~new_n198_ | new_n199_) & ((~new_n200_ & new_n209_) | (~new_n203_ & (new_n200_ | ~new_n209_) & (~new_n200_ | new_n209_))))));
  assign new_n286_ = ((~new_n244_ ^ new_n245_) | (~new_n246_ & new_n247_) | (~new_n248_ & (new_n246_ | ~new_n247_) & (~new_n246_ | new_n247_))) & ((~new_n244_ & new_n245_) | (new_n244_ & ~new_n245_) | ((new_n246_ | ~new_n247_) & (new_n248_ | (~new_n246_ & new_n247_) | (new_n246_ & ~new_n247_)))) & (new_n248_ ^ (~new_n246_ ^ new_n247_)) & ~new_n287_ & ~new_n288_ & new_n289_;
  assign new_n287_ = (new_n251_ ^ (~\a[2]  ^ (new_n250_ & (~new_n47_ | ~new_n249_)))) ^ ((~new_n252_ & new_n253_) | (~new_n254_ & (new_n252_ | ~new_n253_) & (~new_n252_ | new_n253_)));
  assign new_n288_ = ~new_n254_ ^ (~new_n252_ ^ new_n253_);
  assign new_n289_ = ~new_n290_ & (~new_n291_ | ~new_n292_ | ~new_n293_) & (~new_n294_ | ~new_n295_) & \a[0]  & \b[0] ;
  assign new_n290_ = ((\b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] )) ^ (~\a[2]  ^ ((((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] )))) ? ((\b[2]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[1]  & ~\a[0]  & \a[1] ) | (\b[0]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | ((~\b[2]  ^ (\b[0]  | ~\b[1] )) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[0]  & ~\a[0]  & \a[1] ) | (\b[1]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | ((\b[0]  ^ \b[1] ) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | ~\a[2]  | (\a[0]  & \b[0] )) : ((\a[2]  & (~\a[0]  | ~\b[0]  | ((~\b[1]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & ((~\b[0]  ^ \b[1] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))))) | (((~\b[2]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[1]  | \a[0]  | ~\a[1] ) & (~\b[0]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & ((\b[2]  ^ (\b[0]  | ~\b[1] )) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))) ? ((\b[0]  & ~\a[0]  & \a[1] ) | (\b[1]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | ((\b[0]  ^ \b[1] ) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] ))) : ~\a[2] ));
  assign new_n291_ = ~\a[1]  & ~\a[2]  & ~\a[3]  & ~\a[4]  & ~\a[7]  & ~\a[8] ;
  assign new_n292_ = ~\a[13]  & ~\a[14]  & ~\a[11]  & ~\a[12] ;
  assign new_n293_ = ~\a[9]  & ~\a[10]  & ~\a[5]  & ~\a[6]  & ~\a[15]  & ~\a[16]  & ~\a[17]  & ~\a[18] ;
  assign new_n294_ = ~\b[9]  & ~\b[1]  & ~\b[2] ;
  assign new_n295_ = ~\b[7]  & ~\b[8]  & ~\b[5]  & ~\b[6]  & ~\b[3]  & ~\b[4] ;
endmodule


