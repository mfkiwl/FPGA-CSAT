// Benchmark "multiplier_4349_sat" written by ABC on Fri Nov 11 15:24:55 2022

module multiplier_4349_sat ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] ,
    sat  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] ;
  output sat;
  wire new_n23_, new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_,
    new_n30_, new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_,
    new_n37_, new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_,
    new_n44_, new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_,
    new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_,
    new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_,
    new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_,
    new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_,
    new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_,
    new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_,
    new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_,
    new_n100_, new_n101_, new_n102_, new_n103_, new_n104_, new_n105_,
    new_n106_, new_n107_, new_n108_, new_n109_, new_n110_, new_n111_,
    new_n112_, new_n113_, new_n114_, new_n115_, new_n116_, new_n117_,
    new_n118_, new_n119_, new_n120_, new_n121_;
  assign sat = (((~new_n23_ | ~\a[2] ) & ((new_n23_ & \a[2] ) | (~new_n23_ & ~\a[2] ) | ((~new_n77_ | ~\a[2] ) & (new_n78_ | (new_n77_ & \a[2] ) | (~new_n77_ & ~\a[2] ))))) ^ (~new_n101_ ^ (~new_n121_ ^ \a[2] ))) & ((~new_n23_ ^ \a[2] ) ^ ((new_n77_ & \a[2] ) | (~new_n78_ & (~new_n77_ | ~\a[2] ) & (new_n77_ | \a[2] )))) & new_n103_ & (new_n78_ ^ (new_n77_ ^ \a[2] ));
  assign new_n23_ = ((\a[5]  & (new_n67_ | (new_n70_ & \a[8] ) | (~new_n70_ & ~\a[8] )) & (~new_n67_ | (new_n70_ ^ \a[8] ))) | (((new_n73_ & \a[5] ) | (~new_n24_ & (~new_n73_ | ~\a[5] ) & (new_n73_ | \a[5] ))) & (~\a[5]  | (~new_n67_ & (~new_n70_ | ~\a[8] ) & (new_n70_ | \a[8] )) | (new_n67_ & (~new_n70_ ^ \a[8] ))) & (\a[5]  | (~new_n67_ ^ (new_n70_ ^ \a[8] ))))) ^ (\a[5]  ^ (new_n74_ ^ ((new_n70_ & \a[8] ) | (~new_n67_ & (~new_n70_ | ~\a[8] ) & (new_n70_ | \a[8] )))));
  assign new_n24_ = (~new_n25_ | ~\a[5] ) & (new_n49_ | (new_n25_ & \a[5] ) | (~new_n25_ & ~\a[5] ));
  assign new_n25_ = ~new_n26_ ^ (~new_n48_ ^ (~new_n47_ ^ (~new_n46_ ^ (\a[11]  & ~\b[2] ))));
  assign new_n26_ = (~new_n27_ | new_n31_) & (((new_n33_ | ~new_n44_) & (((new_n35_ | ~new_n45_) & (new_n37_ | (~new_n35_ & new_n45_) | (new_n35_ & ~new_n45_))) | (~new_n33_ & new_n44_) | (new_n33_ & ~new_n44_))) | (new_n27_ & ~new_n31_) | (~new_n27_ & new_n31_));
  assign new_n27_ = ~new_n28_ ^ ((\a[11]  & ~\b[1] ) ^ (~new_n30_ | (new_n29_ & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] ))));
  assign new_n28_ = (~\a[11]  | ~\b[0]  | (\b[0]  & (\a[8]  ^ ~\a[9] ) & (\a[9]  | \a[10] ) & (~\a[9]  | ~\a[10] )) | (\b[1]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  ^ ~\a[11] )) | ((\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] )) | (\b[0]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] )) | ((\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] ) & (\b[2]  | ~\b[0]  | ~\b[1] ) & (\b[1]  | \b[2] ) & (~\b[2]  | \b[0]  | ~\b[1] )) | (\b[0]  & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] ) & (\a[8]  ^ ~\a[9] ) & (\a[9]  ^ ~\a[10] )) | (\b[1]  & (\a[8]  ^ ~\a[9] ) & (\a[9]  | \a[10] ) & (~\a[9]  | ~\a[10] )) | (\b[2]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  ^ ~\a[11] ))) & ((\a[11]  ^ (((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  ^ ~\a[10] )) & (~\b[2]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[3]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )))) | (\a[11]  & \b[0]  & (~\b[0]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\b[2]  & \b[0]  & \b[1] ) | (~\b[1]  & ~\b[2] ) | (\b[2]  & ~\b[0]  & \b[1] )) & (~\b[0]  | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  ^ ~\a[10] )) & (~\b[1]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[2]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] ))) | ((~\a[11]  | ~\b[0] ) & ((\b[0]  & (\a[8]  ^ ~\a[9] ) & (\a[9]  | \a[10] ) & (~\a[9]  | ~\a[10] )) | (\b[1]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  ^ ~\a[11] )) | ((\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] )) | ~\a[11]  | (\b[0]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] )) | ((\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] ) & (\b[2]  | ~\b[0]  | ~\b[1] ) & (\b[1]  | \b[2] ) & (~\b[2]  | \b[0]  | ~\b[1] )) | (\b[0]  & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] ) & (\a[8]  ^ ~\a[9] ) & (\a[9]  ^ ~\a[10] )) | (\b[1]  & (\a[8]  ^ ~\a[9] ) & (\a[9]  | \a[10] ) & (~\a[9]  | ~\a[10] )) | (\b[2]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  ^ ~\a[11] )))));
  assign new_n29_ = (\b[3]  ^ \b[4] ) ^ ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] )));
  assign new_n30_ = (~\b[2]  | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  ^ ~\a[10] )) & (~\b[3]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[4]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] ));
  assign new_n31_ = \a[8]  ^ (((new_n32_ ^ \b[6] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[5]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[6]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )));
  assign new_n32_ = (~\b[5]  | ~\b[6] ) & ((~\b[5]  & ~\b[6] ) | (\b[5]  & \b[6] ) | ((~\b[4]  | ~\b[5] ) & ((\b[4]  & \b[5] ) | (~\b[4]  & ~\b[5] ) | ((~\b[3]  | ~\b[4] ) & ((\b[3]  & \b[4] ) | (~\b[3]  & ~\b[4] ) | ((~\b[2]  | ~\b[3] ) & ((~\b[2]  & ~\b[3] ) | (\b[2]  & \b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] ))))))));
  assign new_n33_ = \a[8]  ^ ((~new_n34_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[4]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[5]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[6]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )));
  assign new_n34_ = (~\b[5]  ^ ~\b[6] ) ^ ((\b[4]  & \b[5] ) | ((~\b[4]  | ~\b[5] ) & (\b[4]  | \b[5] ) & ((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] )))))));
  assign new_n35_ = \a[8]  ^ ((~new_n36_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[3]  | (~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[4]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[5]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )));
  assign new_n36_ = (\b[4]  ^ \b[5] ) ^ ((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] )))));
  assign new_n37_ = (~new_n40_ | (\a[8]  ^ (new_n39_ & (~new_n29_ | ~new_n38_)))) & ((~new_n41_ & (new_n42_ | ~new_n43_)) | (new_n40_ & (~\a[8]  ^ (new_n39_ & (~new_n29_ | ~new_n38_)))) | (~new_n40_ & (~\a[8]  | ~new_n39_ | (new_n29_ & new_n38_)) & (\a[8]  | (new_n39_ & (~new_n29_ | ~new_n38_)))));
  assign new_n38_ = (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] );
  assign new_n39_ = (~\b[3]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[4]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[2]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ));
  assign new_n40_ = ((\b[0]  & (\a[8]  ^ ~\a[9] ) & (\a[9]  | \a[10] ) & (~\a[9]  | ~\a[10] )) | (\b[1]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  ^ ~\a[11] )) | ((\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[11]  & \b[0]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ));
  assign new_n41_ = \b[0]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] ) & (~\b[0]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\b[0]  & ~\b[1] ) | (\b[0]  & \b[1] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\b[2]  & \b[0]  & \b[1] ) | (~\b[1]  & ~\b[2] ) | (~\b[0]  & \b[1]  & \b[2] )) & (~\b[1]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[2]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ));
  assign new_n42_ = \a[8]  ^ (((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[3]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[1]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )));
  assign new_n43_ = (\b[0]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] )) ^ ((~\b[0]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\b[0]  & ~\b[1] ) | (\b[0]  & \b[1] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\b[2]  & \b[0]  & \b[1] ) | (~\b[1]  & ~\b[2] ) | (~\b[0]  & \b[1]  & \b[2] )) & (~\b[1]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[2]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )));
  assign new_n44_ = (~\a[11]  ^ (((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  ^ ~\a[10] )) & (~\b[2]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[3]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )))) ^ ((\a[11]  & \b[0] ) ^ ((~\b[0]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\b[2]  & \b[0]  & \b[1] ) | (~\b[1]  & ~\b[2] ) | (\b[2]  & ~\b[0]  & \b[1] )) & (~\b[0]  | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  ^ ~\a[10] )) & (~\b[1]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[2]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] ))));
  assign new_n45_ = (((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\b[2]  & \b[0]  & \b[1] ) | (~\b[1]  & ~\b[2] ) | (\b[2]  & ~\b[0]  & \b[1] )) & (~\b[0]  | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  ^ ~\a[10] )) & (~\b[1]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[2]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] ))) ^ (~\a[11]  | ((~\b[0]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[1]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  ^ ~\a[11] )) & ((~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ))));
  assign new_n46_ = (~new_n36_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[4]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[5]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[3]  | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  ^ ~\a[10] ));
  assign new_n47_ = (new_n28_ | (\a[11]  & ~\b[1]  & (~new_n30_ | (new_n29_ & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] )))) | ((~\a[11]  | \b[1] ) & new_n30_ & (~new_n29_ | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\a[10]  & ~\a[11] ) | (\a[10]  & \a[11] )))) & (~new_n30_ | (new_n29_ & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] ) & (\a[10]  | \a[11] ) & (~\a[10]  | ~\a[11] )) | ~\a[11]  | ~\b[1] );
  assign new_n48_ = \a[8]  ^ (~\b[6]  | (((~\a[6]  ^ ~\a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )) & (new_n32_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ))));
  assign new_n49_ = (~new_n51_ | ~\a[5] ) & (((~\a[5]  | (new_n50_ & ((~new_n35_ & new_n45_) | (~new_n37_ & (new_n35_ | ~new_n45_) & (~new_n35_ | new_n45_)))) | (~new_n50_ & (new_n35_ | ~new_n45_) & (new_n37_ | (~new_n35_ & new_n45_) | (new_n35_ & ~new_n45_)))) & ((\a[5]  & (~new_n50_ | ((new_n35_ | ~new_n45_) & (new_n37_ | (~new_n35_ & new_n45_) | (new_n35_ & ~new_n45_)))) & (new_n50_ | (~new_n35_ & new_n45_) | (~new_n37_ & (new_n35_ | ~new_n45_) & (~new_n35_ | new_n45_)))) | (~\a[5]  & (~new_n50_ ^ ((~new_n35_ & new_n45_) | (~new_n37_ & (new_n35_ | ~new_n45_) & (~new_n35_ | new_n45_))))) | ((new_n66_ | (~new_n37_ & (new_n35_ | ~new_n45_) & (~new_n35_ | new_n45_)) | (new_n37_ & (new_n35_ ^ new_n45_))) & (new_n52_ | (~new_n66_ & (new_n37_ | (~new_n35_ & new_n45_) | (new_n35_ & ~new_n45_)) & (~new_n37_ | (~new_n35_ ^ new_n45_))) | (new_n66_ & (new_n37_ ^ (~new_n35_ ^ new_n45_))))))) | (new_n51_ & \a[5] ) | (~new_n51_ & ~\a[5] ));
  assign new_n50_ = new_n33_ ^ ~new_n44_;
  assign new_n51_ = ((~new_n33_ & new_n44_) | (((~new_n35_ & new_n45_) | (~new_n37_ & (new_n35_ | ~new_n45_) & (~new_n35_ | new_n45_))) & (new_n33_ | ~new_n44_) & (~new_n33_ | new_n44_))) ^ (new_n27_ ^ ~new_n31_);
  assign new_n52_ = (~new_n53_ | new_n54_) & ((new_n53_ & ~new_n54_) | (~new_n53_ & new_n54_) | ((~new_n55_ | new_n56_) & (((new_n57_ | ~new_n65_) & (new_n58_ | (~new_n57_ & new_n65_) | (new_n57_ & ~new_n65_))) | (new_n55_ & ~new_n56_) | (~new_n55_ & new_n56_))));
  assign new_n53_ = (new_n41_ | (~new_n42_ & new_n43_)) ^ (new_n40_ ^ (~\a[8]  ^ (new_n39_ & (~new_n29_ | ~new_n38_))));
  assign new_n54_ = \a[5]  ^ (((new_n32_ ^ \b[6] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[5]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[6]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )));
  assign new_n55_ = new_n42_ ^ ~new_n43_;
  assign new_n56_ = \a[5]  ^ ((~new_n34_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[4]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[5]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[6]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )));
  assign new_n57_ = \a[5]  ^ ((~new_n36_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[3]  | (~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[4]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[5]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )));
  assign new_n58_ = (~new_n61_ | (\a[5]  ^ (new_n60_ & (~new_n29_ | ~new_n59_)))) & ((~new_n62_ & (new_n63_ | ~new_n64_)) | (new_n61_ & (~\a[5]  ^ (new_n60_ & (~new_n29_ | ~new_n59_)))) | (~new_n61_ & (~\a[5]  | ~new_n60_ | (new_n29_ & new_n59_)) & (\a[5]  | (new_n60_ & (~new_n29_ | ~new_n59_)))));
  assign new_n59_ = (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (\a[4]  | \a[5] ) & (~\a[4]  | ~\a[5] );
  assign new_n60_ = (~\b[3]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[4]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[2]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n61_ = ((\b[0]  & (\a[5]  ^ ~\a[6] ) & (\a[6]  | \a[7] ) & (~\a[6]  | ~\a[7] )) | (\b[1]  & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (\a[7]  ^ ~\a[8] )) | ((\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (\a[7]  | \a[8] ) & (~\a[7]  | ~\a[8] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[8]  & \b[0]  & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ));
  assign new_n62_ = \b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (~\b[0]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\b[0]  & ~\b[1] ) | (\b[0]  & \b[1] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\b[2]  & \b[0]  & \b[1] ) | (~\b[1]  & ~\b[2] ) | (~\b[0]  & \b[1]  & \b[2] )) & (~\b[1]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[2]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ));
  assign new_n63_ = \a[5]  ^ (((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[3]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[1]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )));
  assign new_n64_ = (\b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] )) ^ ((~\b[0]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\b[0]  & ~\b[1] ) | (\b[0]  & \b[1] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\b[2]  & \b[0]  & \b[1] ) | (~\b[1]  & ~\b[2] ) | (~\b[0]  & \b[1]  & \b[2] )) & (~\b[1]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[2]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )));
  assign new_n65_ = (~\a[8]  | ((~\b[0]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[1]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & ((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )))) ^ (((~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] ) | (~\b[2]  & \b[0]  & \b[1] ) | (~\b[1]  & ~\b[2] ) | (\b[2]  & ~\b[0]  & \b[1] )) & (~\b[1]  | (~\a[5]  ^ ~\a[6] ) | (~\a[6]  & ~\a[7] ) | (\a[6]  & \a[7] )) & (~\b[2]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\a[7]  ^ ~\a[8] )) & (~\b[0]  | (~\a[6]  ^ ~\a[7] ) | (~\a[5]  ^ ~\a[6] ) | (~\a[7]  & ~\a[8] ) | (\a[7]  & \a[8] )));
  assign new_n66_ = \a[5]  ^ (~\b[6]  | (((~\a[3]  ^ ~\a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )) & (new_n32_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ))));
  assign new_n67_ = (~\a[8]  | (new_n68_ & ((~new_n47_ & (new_n46_ | ~\a[11]  | \b[2] ) & (~new_n46_ | (\a[11]  & ~\b[2] ))) | (new_n46_ & \a[11]  & \b[2] ))) | (~new_n68_ & (new_n47_ | (~new_n46_ & \a[11]  & ~\b[2] ) | (new_n46_ & (~\a[11]  | \b[2] ))) & (~new_n46_ | ~\a[11]  | ~\b[2] ))) & (((new_n48_ | (~new_n47_ & (new_n46_ | ~\a[11]  | \b[2] ) & (~new_n46_ | (\a[11]  & ~\b[2] ))) | (new_n47_ & (new_n46_ ^ (\a[11]  & ~\b[2] )))) & (new_n26_ | (~new_n48_ & (new_n47_ | (~new_n46_ & \a[11]  & ~\b[2] ) | (new_n46_ & (~\a[11]  | \b[2] ))) & (~new_n47_ | (~new_n46_ ^ (\a[11]  & ~\b[2] )))) | (new_n48_ & (new_n47_ ^ (~new_n46_ ^ (\a[11]  & ~\b[2] )))))) | (\a[8]  & (~new_n68_ | ((new_n47_ | (~new_n46_ & \a[11]  & ~\b[2] ) | (new_n46_ & (~\a[11]  | \b[2] ))) & (~new_n46_ | ~\a[11]  | ~\b[2] ))) & (new_n68_ | (~new_n47_ & (new_n46_ | ~\a[11]  | \b[2] ) & (~new_n46_ | (\a[11]  & ~\b[2] ))) | (new_n46_ & \a[11]  & \b[2] ))) | (~\a[8]  & (~new_n68_ ^ ((~new_n47_ & (new_n46_ | ~\a[11]  | \b[2] ) & (~new_n46_ | (\a[11]  & ~\b[2] ))) | (new_n46_ & \a[11]  & \b[2] )))));
  assign new_n68_ = ~new_n69_ ^ (\a[11]  & ~\b[3] );
  assign new_n69_ = (~new_n34_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[5]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[6]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[4]  | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  ^ ~\a[10] ));
  assign new_n70_ = ~new_n71_ ^ (~new_n72_ ^ (\a[11]  & ~\b[4] ));
  assign new_n71_ = ((~new_n69_ & \a[11]  & ~\b[3] ) | (new_n69_ & (~\a[11]  | \b[3] )) | ((new_n47_ | (~new_n46_ & \a[11]  & ~\b[2] ) | (new_n46_ & (~\a[11]  | \b[2] ))) & (~new_n46_ | ~\a[11]  | ~\b[2] ))) & (~new_n69_ | ~\a[11]  | ~\b[3] );
  assign new_n72_ = ((new_n32_ ^ \b[6] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[6]  | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  & ~\a[10] ) | (\a[9]  & \a[10] )) & (~\b[5]  | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] ) | (~\a[9]  ^ ~\a[10] ));
  assign new_n73_ = ((~new_n48_ & (new_n47_ | (~new_n46_ & \a[11]  & ~\b[2] ) | (new_n46_ & (~\a[11]  | \b[2] ))) & (~new_n47_ | (~new_n46_ ^ (\a[11]  & ~\b[2] )))) | (~new_n26_ & (new_n48_ | (~new_n47_ & (new_n46_ | ~\a[11]  | \b[2] ) & (~new_n46_ | (\a[11]  & ~\b[2] ))) | (new_n47_ & (new_n46_ ^ (\a[11]  & ~\b[2] )))) & (~new_n48_ | (~new_n47_ ^ (~new_n46_ ^ (\a[11]  & ~\b[2] )))))) ^ (\a[8]  ^ (new_n68_ ^ ((~new_n47_ & (new_n46_ | ~\a[11]  | \b[2] ) & (~new_n46_ | (\a[11]  & ~\b[2] ))) | (new_n46_ & \a[11]  & \b[2] ))));
  assign new_n74_ = ~\a[8]  ^ (new_n75_ ^ ((~new_n71_ & (new_n72_ | ~\a[11]  | \b[4] ) & (~new_n72_ | (\a[11]  & ~\b[4] ))) | (new_n72_ & \a[11]  & \b[4] )));
  assign new_n75_ = ~new_n76_ ^ (\a[11]  & ~\b[5] );
  assign new_n76_ = \b[6]  & (((~\a[10]  | ~\a[11] ) & (\a[10]  | \a[11] ) & (\a[8]  ^ ~\a[9] ) & (\a[9]  ^ ~\a[10] )) | (~new_n32_ & (~\a[10]  | ~\a[11] ) & (\a[10]  | \a[11] ) & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] )));
  assign new_n77_ = ((new_n73_ & \a[5] ) | (~new_n24_ & (~new_n73_ | ~\a[5] ) & (new_n73_ | \a[5] ))) ^ (\a[5]  ^ (~new_n67_ ^ (new_n70_ ^ \a[8] )));
  assign new_n78_ = (~\a[2]  | (~new_n24_ & (~new_n73_ | ~\a[5] ) & (new_n73_ | \a[5] )) | (new_n24_ & (~new_n73_ ^ \a[5] ))) & (new_n79_ | (\a[2]  & (new_n24_ | (new_n73_ & \a[5] ) | (~new_n73_ & ~\a[5] )) & (~new_n24_ | (new_n73_ ^ \a[5] ))) | (~\a[2]  & (new_n24_ ^ (new_n73_ ^ \a[5] ))));
  assign new_n79_ = (~\a[2]  | (((new_n51_ & \a[5] ) | (~new_n80_ & (~new_n51_ | ~\a[5] ) & (new_n51_ | \a[5] ))) & (~new_n25_ | ~\a[5] ) & (new_n25_ | \a[5] )) | ((~new_n51_ | ~\a[5] ) & (new_n80_ | (new_n51_ & \a[5] ) | (~new_n51_ & ~\a[5] )) & (~new_n25_ ^ \a[5] ))) & (((~\a[2]  | (~new_n80_ & (~new_n51_ | ~\a[5] ) & (new_n51_ | \a[5] )) | (new_n80_ & (~new_n51_ ^ \a[5] ))) & (((~new_n81_ | ~\a[2] ) & ((new_n81_ & \a[2] ) | (~new_n81_ & ~\a[2] ) | ((~new_n82_ | ~\a[2] ) & (new_n83_ | (new_n82_ & \a[2] ) | (~new_n82_ & ~\a[2] ))))) | (\a[2]  & (new_n80_ | (new_n51_ & \a[5] ) | (~new_n51_ & ~\a[5] )) & (~new_n80_ | (new_n51_ ^ \a[5] ))) | (~\a[2]  & (new_n80_ ^ (new_n51_ ^ \a[5] ))))) | (\a[2]  & (((~new_n51_ | ~\a[5] ) & (new_n80_ | (new_n51_ & \a[5] ) | (~new_n51_ & ~\a[5] ))) | (new_n25_ & \a[5] ) | (~new_n25_ & ~\a[5] )) & ((new_n51_ & \a[5] ) | (~new_n80_ & (~new_n51_ | ~\a[5] ) & (new_n51_ | \a[5] )) | (new_n25_ ^ \a[5] ))) | (~\a[2]  & (((~new_n51_ | ~\a[5] ) & (new_n80_ | (new_n51_ & \a[5] ) | (~new_n51_ & ~\a[5] ))) ^ (new_n25_ ^ \a[5] ))));
  assign new_n80_ = (~\a[5]  | (new_n50_ & ((~new_n35_ & new_n45_) | (~new_n37_ & (new_n35_ | ~new_n45_) & (~new_n35_ | new_n45_)))) | (~new_n50_ & (new_n35_ | ~new_n45_) & (new_n37_ | (~new_n35_ & new_n45_) | (new_n35_ & ~new_n45_)))) & ((\a[5]  & (~new_n50_ | ((new_n35_ | ~new_n45_) & (new_n37_ | (~new_n35_ & new_n45_) | (new_n35_ & ~new_n45_)))) & (new_n50_ | (~new_n35_ & new_n45_) | (~new_n37_ & (new_n35_ | ~new_n45_) & (~new_n35_ | new_n45_)))) | (~\a[5]  & (~new_n50_ ^ ((~new_n35_ & new_n45_) | (~new_n37_ & (new_n35_ | ~new_n45_) & (~new_n35_ | new_n45_))))) | ((new_n66_ | (~new_n37_ & (new_n35_ | ~new_n45_) & (~new_n35_ | new_n45_)) | (new_n37_ & (new_n35_ ^ new_n45_))) & (new_n52_ | (~new_n66_ & (new_n37_ | (~new_n35_ & new_n45_) | (new_n35_ & ~new_n45_)) & (~new_n37_ | (~new_n35_ ^ new_n45_))) | (new_n66_ & (new_n37_ ^ (~new_n35_ ^ new_n45_))))));
  assign new_n81_ = (\a[5]  ^ (new_n50_ ^ ((~new_n35_ & new_n45_) | (~new_n37_ & (new_n35_ | ~new_n45_) & (~new_n35_ | new_n45_))))) ^ ((~new_n66_ & (new_n37_ | (~new_n35_ & new_n45_) | (new_n35_ & ~new_n45_)) & (~new_n37_ | (~new_n35_ ^ new_n45_))) | (~new_n52_ & (new_n66_ | (~new_n37_ & (new_n35_ | ~new_n45_) & (~new_n35_ | new_n45_)) | (new_n37_ & (new_n35_ ^ new_n45_))) & (~new_n66_ | (~new_n37_ ^ (~new_n35_ ^ new_n45_)))));
  assign new_n82_ = ~new_n52_ ^ (~new_n66_ ^ (~new_n37_ ^ (~new_n35_ ^ new_n45_)));
  assign new_n83_ = (~new_n85_ | ~\a[2] ) & (((~\a[2]  | (new_n84_ & ((~new_n57_ & new_n65_) | (~new_n58_ & (new_n57_ | ~new_n65_) & (~new_n57_ | new_n65_)))) | (~new_n84_ & (new_n57_ | ~new_n65_) & (new_n58_ | (~new_n57_ & new_n65_) | (new_n57_ & ~new_n65_)))) & ((\a[2]  & (~new_n84_ | ((new_n57_ | ~new_n65_) & (new_n58_ | (~new_n57_ & new_n65_) | (new_n57_ & ~new_n65_)))) & (new_n84_ | (~new_n57_ & new_n65_) | (~new_n58_ & (new_n57_ | ~new_n65_) & (~new_n57_ | new_n65_)))) | (~\a[2]  & (~new_n84_ ^ ((~new_n57_ & new_n65_) | (~new_n58_ & (new_n57_ | ~new_n65_) & (~new_n57_ | new_n65_))))) | ((new_n100_ | (~new_n58_ & (new_n57_ | ~new_n65_) & (~new_n57_ | new_n65_)) | (new_n58_ & (new_n57_ ^ new_n65_))) & (new_n86_ | (~new_n100_ & (new_n58_ | (~new_n57_ & new_n65_) | (new_n57_ & ~new_n65_)) & (~new_n58_ | (~new_n57_ ^ new_n65_))) | (new_n100_ & (new_n58_ ^ (~new_n57_ ^ new_n65_))))))) | (new_n85_ & \a[2] ) | (~new_n85_ & ~\a[2] ));
  assign new_n84_ = new_n55_ ^ ~new_n56_;
  assign new_n85_ = (new_n53_ ^ ~new_n54_) ^ ((new_n55_ & ~new_n56_) | (((~new_n57_ & new_n65_) | (~new_n58_ & (new_n57_ | ~new_n65_) & (~new_n57_ | new_n65_))) & (~new_n55_ | new_n56_) & (new_n55_ | ~new_n56_)));
  assign new_n86_ = (new_n87_ | ~new_n88_) & ((new_n87_ & ~new_n88_) | (~new_n87_ & new_n88_) | ((new_n89_ | ~new_n91_) & ((new_n89_ & ~new_n91_) | (~new_n89_ & new_n91_) | (~new_n92_ & (~new_n94_ | new_n95_)))));
  assign new_n87_ = \a[2]  ^ (((~new_n32_ ^ ~\b[6] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[5]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[6]  | \a[0]  | ~\a[1] ));
  assign new_n88_ = (new_n62_ | (~new_n63_ & new_n64_)) ^ (new_n61_ ^ (~\a[5]  ^ (new_n60_ & (~new_n29_ | ~new_n59_))));
  assign new_n89_ = \a[2]  ^ (new_n90_ & (~new_n34_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )));
  assign new_n90_ = (~\b[4]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[6]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[5]  | \a[0]  | ~\a[1] );
  assign new_n91_ = new_n63_ ^ ~new_n64_;
  assign new_n92_ = new_n93_ & (~\a[2]  ^ ((~new_n36_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[3]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | \a[0]  | \a[1] ) & (~\b[5]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[4]  | \a[0]  | ~\a[1] )));
  assign new_n93_ = (~\a[5]  | ((~\b[0]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[1]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & ((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )))) ^ (((~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] ) | (~\b[2]  & \b[0]  & \b[1] ) | (~\b[1]  & ~\b[2] ) | (\b[2]  & ~\b[0]  & \b[1] )) & (~\b[1]  | (~\a[2]  ^ ~\a[3] ) | (~\a[3]  & ~\a[4] ) | (\a[3]  & \a[4] )) & (~\b[2]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\a[4]  ^ ~\a[5] )) & (~\b[0]  | (~\a[3]  ^ ~\a[4] ) | (~\a[2]  ^ ~\a[3] ) | (~\a[4]  & ~\a[5] ) | (\a[4]  & \a[5] )));
  assign new_n94_ = new_n93_ ^ (~\a[2]  ^ ((~new_n36_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[3]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | \a[0]  | \a[1] ) & (~\b[5]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[4]  | \a[0]  | ~\a[1] )));
  assign new_n95_ = (new_n96_ | ~new_n97_) & (new_n98_ | new_n99_ | (new_n96_ & ~new_n97_));
  assign new_n96_ = \a[2]  ^ ((((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((\b[2]  | \b[3] ) & (~\b[2]  | ~\b[3] ) & \b[1]  & (\b[0]  | \b[2] )))) | ((~\b[3]  ^ \b[4] ) & (~\b[2]  | ~\b[3] ) & ((~\b[2]  & ~\b[3] ) | (\b[2]  & \b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[2]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[4]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[3]  | \a[0]  | ~\a[1] ));
  assign new_n97_ = ((\b[0]  & (\a[2]  ^ ~\a[3] ) & (\a[3]  | \a[4] ) & (~\a[3]  | ~\a[4] )) | (\b[1]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (\a[4]  ^ ~\a[5] )) | ((\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (\a[4]  | \a[5] ) & (~\a[4]  | ~\a[5] ) & (~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ))) ^ (\a[5]  & \b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ));
  assign new_n98_ = (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (\a[2]  ^ ((~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] ) & (((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))))) & (~\a[2]  | (\a[0]  & \b[0] ) | (\b[1]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[0]  & ~\a[0]  & \a[1] ) | ((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | ((\b[2]  | ~\b[0]  | ~\b[1] ) & (\b[1]  | \b[2] ) & (~\b[2]  | \b[0]  | ~\b[1] ) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[0]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[2]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[1]  & ~\a[0]  & \a[1] ));
  assign new_n99_ = (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\a[2]  | (\b[1]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[3]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[2]  & ~\a[0]  & \a[1] ) | (((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )) & ((\b[2]  ^ \b[3] ) | (\b[1]  & (\b[0]  | \b[2] ))) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] ))) & (\a[2]  | ((~\b[1]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[3]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[2]  | \a[0]  | ~\a[1] ) & (((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))));
  assign new_n100_ = \a[2]  ^ (~\b[6]  | ((\a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (new_n32_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))));
  assign new_n101_ = ((~\a[5]  | (new_n74_ & ((new_n70_ & \a[8] ) | (~new_n67_ & (~new_n70_ | ~\a[8] ) & (new_n70_ | \a[8] )))) | (~new_n74_ & (~new_n70_ | ~\a[8] ) & (new_n67_ | (new_n70_ & \a[8] ) | (~new_n70_ & ~\a[8] )))) & (((~\a[5]  | (~new_n67_ & (~new_n70_ | ~\a[8] ) & (new_n70_ | \a[8] )) | (new_n67_ & (~new_n70_ ^ \a[8] ))) & (((~new_n73_ | ~\a[5] ) & (new_n24_ | (new_n73_ & \a[5] ) | (~new_n73_ & ~\a[5] ))) | (\a[5]  & (new_n67_ | (new_n70_ & \a[8] ) | (~new_n70_ & ~\a[8] )) & (~new_n67_ | (new_n70_ ^ \a[8] ))) | (~\a[5]  & (new_n67_ ^ (new_n70_ ^ \a[8] ))))) | (\a[5]  & (~new_n74_ | ((~new_n70_ | ~\a[8] ) & (new_n67_ | (new_n70_ & \a[8] ) | (~new_n70_ & ~\a[8] )))) & (new_n74_ | (new_n70_ & \a[8] ) | (~new_n67_ & (~new_n70_ | ~\a[8] ) & (new_n70_ | \a[8] )))) | (~\a[5]  & (~new_n74_ ^ ((new_n70_ & \a[8] ) | (~new_n67_ & (~new_n70_ | ~\a[8] ) & (new_n70_ | \a[8] ))))))) ^ (~new_n102_ ^ (\a[5]  ^ ~\a[8] ));
  assign new_n102_ = ((~new_n76_ ^ (\a[11]  & ~\b[5] )) | ((~new_n72_ | ~\a[11]  | ~\b[4] ) & (new_n71_ | (~new_n72_ & \a[11]  & ~\b[4] ) | (new_n72_ & (~\a[11]  | \b[4] ))))) & (new_n76_ | ~\a[11]  | ~\b[5] );
  assign new_n103_ = ~new_n104_ & new_n105_ & (new_n79_ ^ (\a[2]  ^ (~new_n24_ ^ (~new_n73_ ^ ~\a[5] ))));
  assign new_n104_ = ((\a[2]  & (new_n80_ | (new_n51_ & \a[5] ) | (~new_n51_ & ~\a[5] )) & (~new_n80_ | (new_n51_ ^ \a[5] ))) | (((new_n81_ & \a[2] ) | ((~new_n81_ | ~\a[2] ) & (new_n81_ | \a[2] ) & ((new_n82_ & \a[2] ) | (~new_n83_ & (~new_n82_ | ~\a[2] ) & (new_n82_ | \a[2] ))))) & (~\a[2]  | (~new_n80_ & (~new_n51_ | ~\a[5] ) & (new_n51_ | \a[5] )) | (new_n80_ & (~new_n51_ ^ \a[5] ))) & (\a[2]  | (~new_n80_ ^ (new_n51_ ^ \a[5] ))))) ^ (\a[2]  ^ (((new_n51_ & \a[5] ) | (~new_n80_ & (~new_n51_ | ~\a[5] ) & (new_n51_ | \a[5] ))) ^ (new_n25_ ^ \a[5] )));
  assign new_n105_ = ((~new_n106_ ^ \a[2] ) ^ ((new_n81_ & \a[2] ) | ((~new_n81_ | ~\a[2] ) & (new_n81_ | \a[2] ) & ((new_n82_ & \a[2] ) | ((~new_n82_ | ~\a[2] ) & (new_n82_ | \a[2] ) & ((new_n85_ & \a[2] ) | (~new_n107_ & (new_n85_ | \a[2] ) & (~new_n85_ | ~\a[2] )))))))) & ((new_n81_ ^ \a[2] ) | (new_n82_ & \a[2] ) | ((~new_n82_ | ~\a[2] ) & (new_n82_ | \a[2] ) & ((new_n85_ & \a[2] ) | (~new_n107_ & (new_n85_ | \a[2] ) & (~new_n85_ | ~\a[2] ))))) & ((new_n81_ & \a[2] ) | (~new_n81_ & ~\a[2] ) | ((~new_n82_ | ~\a[2] ) & ((new_n82_ & \a[2] ) | (~new_n82_ & ~\a[2] ) | ((~new_n85_ | ~\a[2] ) & (new_n107_ | (~new_n85_ & ~\a[2] ) | (new_n85_ & \a[2] )))))) & ((~new_n82_ ^ \a[2] ) ^ ((new_n85_ & \a[2] ) | (~new_n107_ & (new_n85_ | \a[2] ) & (~new_n85_ | ~\a[2] )))) & new_n108_ & (new_n107_ ^ (~new_n85_ ^ ~\a[2] ));
  assign new_n106_ = ((\a[5]  & (~new_n50_ | ((new_n35_ | ~new_n45_) & (new_n37_ | (~new_n35_ & new_n45_) | (new_n35_ & ~new_n45_)))) & (new_n50_ | (~new_n35_ & new_n45_) | (~new_n37_ & (new_n35_ | ~new_n45_) & (~new_n35_ | new_n45_)))) | ((~\a[5]  | (new_n50_ & ((~new_n35_ & new_n45_) | (~new_n37_ & (new_n35_ | ~new_n45_) & (~new_n35_ | new_n45_)))) | (~new_n50_ & (new_n35_ | ~new_n45_) & (new_n37_ | (~new_n35_ & new_n45_) | (new_n35_ & ~new_n45_)))) & (\a[5]  | (new_n50_ ^ ((~new_n35_ & new_n45_) | (~new_n37_ & (new_n35_ | ~new_n45_) & (~new_n35_ | new_n45_))))) & ((~new_n66_ & (new_n37_ | (~new_n35_ & new_n45_) | (new_n35_ & ~new_n45_)) & (~new_n37_ | (~new_n35_ ^ new_n45_))) | (~new_n52_ & (new_n66_ | (~new_n37_ & (new_n35_ | ~new_n45_) & (~new_n35_ | new_n45_)) | (new_n37_ & (new_n35_ ^ new_n45_))) & (~new_n66_ | (~new_n37_ ^ (~new_n35_ ^ new_n45_))))))) ^ (new_n51_ ^ \a[5] );
  assign new_n107_ = (~\a[2]  | (((~new_n57_ & new_n65_) | (~new_n58_ & (new_n57_ | ~new_n65_) & (~new_n57_ | new_n65_))) & (~new_n55_ | new_n56_) & (new_n55_ | ~new_n56_)) | ((new_n57_ | ~new_n65_) & (new_n58_ | (~new_n57_ & new_n65_) | (new_n57_ & ~new_n65_)) & (~new_n55_ ^ ~new_n56_))) & (((new_n100_ | (~new_n58_ & (new_n57_ | ~new_n65_) & (~new_n57_ | new_n65_)) | (new_n58_ & (new_n57_ ^ new_n65_))) & (new_n86_ | (~new_n100_ & (new_n58_ | (~new_n57_ & new_n65_) | (new_n57_ & ~new_n65_)) & (~new_n58_ | (~new_n57_ ^ new_n65_))) | (new_n100_ & (new_n58_ ^ (~new_n57_ ^ new_n65_))))) | (\a[2]  & (((new_n57_ | ~new_n65_) & (new_n58_ | (~new_n57_ & new_n65_) | (new_n57_ & ~new_n65_))) | (new_n55_ & ~new_n56_) | (~new_n55_ & new_n56_)) & ((~new_n57_ & new_n65_) | (~new_n58_ & (new_n57_ | ~new_n65_) & (~new_n57_ | new_n65_)) | (new_n55_ ^ ~new_n56_))) | (~\a[2]  & (((new_n57_ | ~new_n65_) & (new_n58_ | (~new_n57_ & new_n65_) | (new_n57_ & ~new_n65_))) ^ (new_n55_ ^ ~new_n56_))));
  assign new_n108_ = (~new_n112_ ^ (new_n109_ | (~new_n109_ & ~new_n111_ & ((~new_n87_ & new_n88_) | (~new_n110_ & (new_n87_ | ~new_n88_) & (~new_n87_ | new_n88_)))))) & ((new_n109_ | new_n111_) ^ ((~new_n87_ & new_n88_) | (~new_n110_ & (new_n87_ | ~new_n88_) & (~new_n87_ | new_n88_)))) & (~new_n110_ | (~new_n87_ ^ new_n88_)) & new_n113_ & (new_n110_ | (~new_n87_ & new_n88_) | (new_n87_ & ~new_n88_));
  assign new_n109_ = ~new_n100_ & (new_n58_ | (~new_n57_ & new_n65_) | (new_n57_ & ~new_n65_)) & (~new_n58_ | (~new_n57_ ^ new_n65_));
  assign new_n110_ = (new_n89_ | ~new_n91_) & ((new_n89_ & ~new_n91_) | (~new_n89_ & new_n91_) | (~new_n92_ & (~new_n94_ | new_n95_)));
  assign new_n111_ = new_n100_ & (new_n58_ ^ (~new_n57_ ^ new_n65_));
  assign new_n112_ = \a[2]  ^ ((new_n55_ ^ ~new_n56_) ^ ((~new_n57_ & new_n65_) | (~new_n58_ & (new_n57_ | ~new_n65_) & (~new_n57_ | new_n65_))));
  assign new_n113_ = (new_n114_ | new_n92_ | (new_n94_ & ((~new_n96_ & new_n97_) | (~new_n98_ & (~new_n96_ | new_n97_) & ~new_n99_)))) & (~new_n114_ | (~new_n92_ & (~new_n94_ | ((new_n96_ | ~new_n97_) & (new_n98_ | (new_n96_ & ~new_n97_) | new_n99_))))) & (new_n94_ | (~new_n96_ & new_n97_) | (~new_n98_ & (~new_n96_ | new_n97_) & ~new_n99_)) & (~new_n94_ | ((new_n96_ | ~new_n97_) & (new_n98_ | (new_n96_ & ~new_n97_) | new_n99_))) & (new_n96_ | ~new_n97_) & new_n115_ & ~new_n99_ & new_n98_ & (~new_n96_ | new_n97_);
  assign new_n114_ = (new_n63_ ^ ~new_n64_) ^ (~\a[2]  ^ (new_n90_ & (~new_n34_ | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ))));
  assign new_n115_ = ~new_n116_ & ~new_n117_ & ~new_n118_ & new_n120_ & (~new_n119_ | \a[11]  | \a[7]  | \a[8] );
  assign new_n116_ = (~\a[2]  | (\a[0]  & \b[0] )) & ((\b[0]  & \b[1] ) | (~\b[0]  & ~\b[1] ) | ~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[1]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[0]  | \a[0]  | ~\a[1] ) & (~\b[0]  | \a[0]  | \a[1]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] )) & (~\b[2]  | ~\a[0]  | (~\a[1]  ^ ~\a[2] )) & (~\b[1]  | \a[0]  | ~\a[1] ) & (~\a[0]  | (~\a[1]  & ~\a[2] ) | (\a[1]  & \a[2] ) | (~\b[2]  & \b[0]  & \b[1] ) | (~\b[1]  & ~\b[2] ) | (\b[2]  & ~\b[0]  & \b[1] ));
  assign new_n117_ = ((\b[0]  & ~\a[0]  & ~\a[1]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[2]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[1]  & ~\a[0]  & \a[1] ) | (\a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] ) & (\b[2]  | ~\b[0]  | ~\b[1] ) & (\b[1]  | \b[2] ) & (~\b[2]  | \b[0]  | ~\b[1] ))) & \a[2]  & \a[0]  & \b[0] ;
  assign new_n118_ = (((~\b[0]  | ~\b[1] ) & (\b[0]  | \b[1] ) & \a[0]  & (\a[1]  | \a[2] ) & (~\a[1]  | ~\a[2] )) | (\b[1]  & \a[0]  & (\a[1]  ^ ~\a[2] )) | (\b[0]  & ~\a[0]  & \a[1] )) & (~\a[2]  | ~\a[0]  | ~\b[0] );
  assign new_n119_ = ~\a[5]  & ~\a[6]  & ~\a[9]  & ~\a[10]  & ~\a[1]  & ~\a[2]  & ~\a[3]  & ~\a[4] ;
  assign new_n120_ = \a[0]  & \b[0]  & (\b[1]  | \b[2]  | \b[3]  | \b[4]  | \b[5]  | \b[6] );
  assign new_n121_ = ((~\a[8]  | (~new_n75_ & ((~new_n71_ & (new_n72_ | ~\a[11]  | \b[4] ) & (~new_n72_ | (\a[11]  & ~\b[4] ))) | (new_n72_ & \a[11]  & \b[4] ))) | (new_n75_ & (new_n71_ | (~new_n72_ & \a[11]  & ~\b[4] ) | (new_n72_ & (~\a[11]  | \b[4] ))) & (~new_n72_ | ~\a[11]  | ~\b[4] ))) & (((~\a[8]  | (~new_n71_ & (new_n72_ | ~\a[11]  | \b[4] ) & (~new_n72_ | (\a[11]  & ~\b[4] ))) | (new_n71_ & (new_n72_ ^ (\a[11]  & ~\b[4] )))) & (new_n67_ | (\a[8]  & (new_n71_ | (~new_n72_ & \a[11]  & ~\b[4] ) | (new_n72_ & (~\a[11]  | \b[4] ))) & (~new_n71_ | (~new_n72_ ^ (\a[11]  & ~\b[4] )))) | (~\a[8]  & (new_n71_ ^ (~new_n72_ ^ (\a[11]  & ~\b[4] )))))) | (\a[8]  & (new_n75_ | ((new_n71_ | (~new_n72_ & \a[11]  & ~\b[4] ) | (new_n72_ & (~\a[11]  | \b[4] ))) & (~new_n72_ | ~\a[11]  | ~\b[4] ))) & (~new_n75_ | (~new_n71_ & (new_n72_ | ~\a[11]  | \b[4] ) & (~new_n72_ | (\a[11]  & ~\b[4] ))) | (new_n72_ & \a[11]  & \b[4] ))) | (~\a[8]  & (new_n75_ ^ ((~new_n71_ & (new_n72_ | ~\a[11]  | \b[4] ) & (~new_n72_ | (\a[11]  & ~\b[4] ))) | (new_n72_ & \a[11]  & \b[4] )))))) ^ (~\a[11]  | \b[6] );
endmodule


