// Benchmark "multiplier_248521_sat" written by ABC on Tue Jan 10 14:28:03 2023

module multiplier_248521_sat ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    sat  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] ,
    \b[7] , \b[8] ;
  output sat;
  wire new_n30_, new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_,
    new_n37_, new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_,
    new_n44_, new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_,
    new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_,
    new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_,
    new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_,
    new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_,
    new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_,
    new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_,
    new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_,
    new_n100_, new_n101_, new_n102_, new_n103_, new_n104_, new_n105_,
    new_n106_, new_n107_, new_n108_, new_n109_, new_n110_, new_n111_,
    new_n112_, new_n113_, new_n114_, new_n115_, new_n116_, new_n117_,
    new_n118_, new_n119_, new_n120_, new_n121_, new_n122_, new_n123_,
    new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_,
    new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_,
    new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_,
    new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_,
    new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_,
    new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_,
    new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_,
    new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_,
    new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_;
  assign sat = (((new_n30_ & \a[2] ) | ((~new_n30_ | ~\a[2] ) & (new_n30_ | \a[2] ) & ((new_n160_ & \a[2] ) | (~new_n162_ & (~new_n160_ | ~\a[2] ) & (new_n160_ | \a[2] ))))) ^ (new_n221_ ^ (~new_n198_ ^ ~new_n222_))) & new_n199_ & ((~new_n30_ ^ \a[2] ) ^ ((new_n160_ & \a[2] ) | (~new_n162_ & (~new_n160_ | ~\a[2] ) & (new_n160_ | \a[2] ))));
  assign new_n30_ = ((new_n152_ & \a[5] ) | (~new_n31_ & (~new_n152_ | ~\a[5] ) & (new_n152_ | \a[5] ))) ^ (\a[5]  ^ (~new_n156_ ^ (~\a[8]  ^ (~new_n157_ ^ (~new_n158_ ^ \a[11] )))));
  assign new_n31_ = (~new_n32_ | ~\a[5] ) & ((new_n32_ & \a[5] ) | (~new_n32_ & ~\a[5] ) | ((~new_n118_ | ~\a[5] ) & (new_n119_ | (new_n118_ & \a[5] ) | (~new_n118_ & ~\a[5] ))));
  assign new_n32_ = ((\a[8]  & ((~new_n116_ & ~\a[11] ) | (new_n116_ & \a[11] ) | ((~new_n91_ | ~\a[11] ) & (new_n117_ | (new_n91_ & \a[11] ) | (~new_n91_ & ~\a[11] )))) & ((~new_n116_ ^ ~\a[11] ) | (new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] )))) | (~new_n65_ & (~\a[8]  | ((new_n116_ | \a[11] ) & (~new_n116_ | ~\a[11] ) & ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] )))) | ((new_n116_ ^ ~\a[11] ) & (~new_n91_ | ~\a[11] ) & (new_n117_ | (new_n91_ & \a[11] ) | (~new_n91_ & ~\a[11] )))) & (\a[8]  | ((~new_n116_ ^ ~\a[11] ) ^ ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] ))))))) ^ (\a[8]  ^ (((new_n116_ & \a[11] ) | ((new_n116_ | \a[11] ) & (~new_n116_ | ~\a[11] ) & ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] ))))) ^ (~new_n33_ ^ ~\a[11] )));
  assign new_n33_ = ~new_n34_ ^ (~new_n61_ & (~new_n63_ | (~new_n39_ & ~new_n64_)));
  assign new_n34_ = (new_n35_ ^ \a[14] ) ^ ((new_n38_ & \a[16]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) | (\b[7]  & ~\a[16]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) | (\b[5]  & (~\a[14]  ^ \a[15] ) & \a[15]  & \a[16] ) | (\b[6]  & (~\a[14]  ^ \a[15] ) & (~\a[15]  | ~\a[16] ) & (\a[15]  | \a[16] )));
  assign new_n35_ = \b[8]  & (((~\a[13]  | ~\a[14] ) & (\a[13]  | \a[14] ) & (~\a[12]  ^ \a[13] ) & (~\a[11]  ^ \a[12] )) | (~new_n36_ & (~\a[13]  | ~\a[14] ) & (\a[13]  | \a[14] ) & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] )));
  assign new_n36_ = (~\b[7]  | ~\b[8] ) & (new_n37_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ));
  assign new_n37_ = (~\b[6]  | ~\b[7] ) & (((~\b[5]  | ~\b[6] ) & (((~\b[4]  | ~\b[5] ) & (((~\b[3]  | ~\b[4] ) & ((\b[3]  & \b[4] ) | (~\b[3]  & ~\b[4] ) | ((~\b[2]  | ~\b[3] ) & ((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] ))))) | (\b[4]  & \b[5] ) | (~\b[4]  & ~\b[5] ))) | (\b[5]  & \b[6] ) | (~\b[5]  & ~\b[6] ))) | (\b[6]  & \b[7] ) | (~\b[6]  & ~\b[7] ));
  assign new_n38_ = ((\b[5]  & \b[6] ) | (((\b[4]  & \b[5] ) | (((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))) & (~\b[4]  | ~\b[5] ) & (\b[4]  | \b[5] ))) & (~\b[5]  | ~\b[6] ) & (\b[5]  | \b[6] ))) ^ (\b[6]  ^ \b[7] );
  assign new_n39_ = new_n54_ & ((~new_n40_ & ~new_n41_) | ((new_n40_ | new_n41_) & (~new_n40_ | ~new_n41_) & ((~new_n43_ & ~new_n59_) | ((new_n43_ | new_n59_) & (~new_n43_ | ~new_n59_) & ((~new_n45_ & ~new_n60_) | (~new_n47_ & (new_n45_ | new_n60_) & (~new_n45_ | ~new_n60_)))))));
  assign new_n40_ = \a[14]  ^ ((~new_n38_ | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] )) & (~\b[5]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[12]  ^ \a[13] ) | (\a[11]  ^ \a[12] )) & (~\b[6]  | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] ) | (\a[11]  ^ \a[12] )) & (~\b[7]  | (\a[13]  ^ \a[14] ) | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] )));
  assign new_n41_ = (~new_n42_ | ~\a[16]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] )) & (~\b[4]  | \a[16]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] )) & (~\b[2]  | ~\a[15]  | ~\a[16]  | (\a[14]  ^ \a[15] )) & (~\b[3]  | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] ) | (\a[14]  ^ \a[15] ));
  assign new_n42_ = (\b[3]  ^ \b[4] ) ^ ((\b[2]  & \b[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )));
  assign new_n43_ = \a[14]  ^ ((~new_n44_ | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] )) & (~\b[4]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[12]  ^ \a[13] ) | (\a[11]  ^ \a[12] )) & (~\b[5]  | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] ) | (\a[11]  ^ \a[12] )) & (~\b[6]  | (\a[13]  ^ \a[14] ) | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] )));
  assign new_n44_ = ((\b[4]  & \b[5] ) | (((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))) & (~\b[4]  | ~\b[5] ) & (\b[4]  | \b[5] ))) ^ (\b[5]  ^ \b[6] );
  assign new_n45_ = \a[14]  ^ ((~new_n46_ | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] )) & (~\b[3]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[12]  ^ \a[13] ) | (\a[11]  ^ \a[12] )) & (~\b[4]  | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] ) | (\a[11]  ^ \a[12] )) & (~\b[5]  | (\a[13]  ^ \a[14] ) | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] )));
  assign new_n46_ = ((\b[3]  & \b[4] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] ))))) ^ (\b[4]  ^ \b[5] );
  assign new_n47_ = (new_n50_ | (\a[14]  ^ (new_n49_ & (~new_n48_ | ~new_n42_)))) & ((~new_n51_ & (new_n52_ | ~new_n53_)) | (~new_n50_ & (~\a[14]  ^ (new_n49_ & (~new_n48_ | ~new_n42_)))) | (new_n50_ & (~\a[14]  | ~new_n49_ | (new_n48_ & new_n42_)) & (\a[14]  | (new_n49_ & (~new_n48_ | ~new_n42_)))));
  assign new_n48_ = (~\a[13]  | ~\a[14] ) & (\a[13]  | \a[14] ) & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] );
  assign new_n49_ = (~\b[2]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[12]  ^ \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[3]  | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[4]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ));
  assign new_n50_ = (~\b[0]  | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[1]  | \a[16]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\a[16]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\b[0]  ^ \b[1] ));
  assign new_n51_ = \b[0]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] ) & (~\b[0]  | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[1]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\b[0]  ^ \b[1] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[0]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[12]  ^ \a[13] ) | (~\a[11]  ^ ~\a[12] )) & ((\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\b[2]  & (\b[0]  | ~\b[1] )) | (\b[2]  & ~\b[0]  & \b[1] )) & (~\b[1]  | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[2]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ));
  assign new_n52_ = \a[14]  ^ (((\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[1]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[12]  ^ \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[2]  | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[3]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )));
  assign new_n53_ = (\b[0]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) ^ ((~\b[0]  | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[1]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\b[0]  ^ \b[1] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & (~\b[0]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[12]  ^ \a[13] ) | (~\a[11]  ^ ~\a[12] )) & ((\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\b[2]  & (\b[0]  | ~\b[1] )) | (\b[2]  & ~\b[0]  & \b[1] )) & (~\b[1]  | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[2]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )));
  assign new_n54_ = (~\a[14]  ^ (new_n56_ & (~new_n48_ | (~new_n37_ & new_n55_) | (new_n37_ & ~new_n55_)))) ^ (~new_n58_ | (new_n57_ & new_n46_));
  assign new_n55_ = ~\b[7]  ^ ~\b[8] ;
  assign new_n56_ = (~\b[6]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[12]  ^ \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[7]  | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[8]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ));
  assign new_n57_ = \a[16]  & (\a[14]  | \a[15] ) & (~\a[14]  | ~\a[15] );
  assign new_n58_ = (~\b[5]  | \a[16]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[3]  | ~\a[15]  | ~\a[16]  | (~\a[14]  ^ ~\a[15] )) & (~\b[4]  | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] ) | (~\a[14]  ^ ~\a[15] ));
  assign new_n59_ = (~\a[16]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[3]  | \a[16]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\b[2]  | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[1]  | ~\a[15]  | ~\a[16]  | (~\a[14]  ^ ~\a[15] ));
  assign new_n60_ = (~\b[0]  | ~\a[15]  | ~\a[16]  | (~\a[14]  ^ ~\a[15] )) & (~\b[1]  | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] ) | (~\a[14]  ^ ~\a[15] )) & (~\b[2]  | \a[16]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] )) & (~\a[16]  | (~\a[14]  & ~\a[15] ) | (\a[14]  & \a[15] ) | (~\b[2]  & (\b[0]  | ~\b[1] )) | (\b[2]  & ~\b[0]  & \b[1] ));
  assign new_n61_ = ((new_n44_ & \a[16]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) | (\b[6]  & ~\a[16]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) | (\b[4]  & (~\a[14]  ^ \a[15] ) & \a[15]  & \a[16] ) | (\b[5]  & (~\a[14]  ^ \a[15] ) & (~\a[15]  | ~\a[16] ) & (\a[15]  | \a[16] ))) & (new_n62_ ^ ~\a[14] );
  assign new_n62_ = ((\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[11]  & \a[12] ) | (~\a[11]  & ~\a[12] ) | (~\b[8]  ^ ((\b[7]  & \b[8] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))))) & (~\b[7]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[12]  ^ \a[13] ) | (\a[11]  ^ \a[12] )) & (~\b[8]  | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] ) | (\a[11]  ^ \a[12] ));
  assign new_n63_ = ((new_n44_ & \a[16]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) | (\b[6]  & ~\a[16]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) | (\b[4]  & (~\a[14]  ^ \a[15] ) & \a[15]  & \a[16] ) | (\b[5]  & (~\a[14]  ^ \a[15] ) & (~\a[15]  | ~\a[16] ) & (\a[15]  | \a[16] ))) ^ (new_n62_ ^ ~\a[14] );
  assign new_n64_ = (~\a[14]  ^ (new_n56_ & (~new_n48_ | (~new_n37_ & new_n55_) | (new_n37_ & ~new_n55_)))) & (~new_n58_ | (new_n57_ & new_n46_));
  assign new_n65_ = (~\a[8]  | (new_n90_ & (new_n66_ | (~new_n69_ & new_n89_))) | (~new_n90_ & ~new_n66_ & (new_n69_ | ~new_n89_))) & (((~\a[8]  | (~new_n69_ & new_n89_) | (new_n69_ & ~new_n89_)) & ((\a[8]  & (new_n69_ | ~new_n89_) & (~new_n69_ | new_n89_)) | (~\a[8]  & (new_n69_ ^ new_n89_)) | ((~new_n92_ | ~\a[8] ) & ((new_n92_ & \a[8] ) | (~new_n92_ & ~\a[8] ) | ((~new_n93_ | ~\a[8] ) & (new_n94_ | (new_n93_ & \a[8] ) | (~new_n93_ & ~\a[8] ))))))) | (\a[8]  & (~new_n90_ | (~new_n66_ & (new_n69_ | ~new_n89_))) & (new_n90_ | new_n66_ | (~new_n69_ & new_n89_))) | (~\a[8]  & (~new_n90_ ^ (new_n66_ | (~new_n69_ & new_n89_)))));
  assign new_n66_ = new_n67_ & ~new_n68_;
  assign new_n67_ = (~new_n40_ ^ ~new_n41_) ^ ((~new_n43_ & ~new_n59_) | (((~new_n45_ & ~new_n60_) | (~new_n47_ & (new_n45_ | new_n60_) & (~new_n45_ | ~new_n60_))) & (new_n43_ | new_n59_) & (~new_n43_ | ~new_n59_)));
  assign new_n68_ = \a[11]  ^ (~\b[8]  | ((new_n36_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] )) & ((\a[9]  ^ \a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\a[8]  ^ \a[9] ))));
  assign new_n69_ = (~new_n70_ | new_n88_) & ((~new_n71_ & (new_n73_ | ~new_n87_)) | (new_n70_ & ~new_n88_) | (~new_n70_ & new_n88_));
  assign new_n70_ = (new_n43_ ^ new_n59_) ^ ((~new_n45_ & ~new_n60_) | (~new_n47_ & (new_n45_ | new_n60_) & (~new_n45_ | ~new_n60_)));
  assign new_n71_ = ~new_n72_ & (new_n47_ | (new_n45_ & new_n60_) | (~new_n45_ & ~new_n60_)) & (~new_n47_ | (new_n45_ ^ new_n60_));
  assign new_n72_ = \a[11]  ^ (((\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n37_ & (~\b[7]  ^ \b[8] ))) & (~\b[7]  | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] ) | (\a[8]  ^ \a[9] )) & (~\b[8]  | (\a[10]  ^ \a[11] ) | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] )) & (~\b[6]  | (\a[9]  ^ \a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\a[8]  ^ \a[9] )));
  assign new_n73_ = (new_n74_ | ~new_n75_) & ((new_n74_ & ~new_n75_) | (~new_n74_ & new_n75_) | ((~new_n76_ | new_n77_) & (((new_n78_ | ~new_n86_) & (new_n79_ | (~new_n78_ & new_n86_) | (new_n78_ & ~new_n86_))) | (~new_n76_ & new_n77_) | (new_n76_ & ~new_n77_))));
  assign new_n74_ = \a[11]  ^ ((~new_n38_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] )) & (~\b[6]  | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] ) | (\a[8]  ^ \a[9] )) & (~\b[7]  | (\a[10]  ^ \a[11] ) | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] )) & (~\b[5]  | (\a[9]  ^ \a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\a[8]  ^ \a[9] )));
  assign new_n75_ = (new_n51_ | (~new_n52_ & new_n53_)) ^ (~new_n50_ ^ (~\a[14]  ^ (new_n49_ & (~new_n48_ | ~new_n42_))));
  assign new_n76_ = new_n52_ ^ ~new_n53_;
  assign new_n77_ = \a[11]  ^ ((~new_n44_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] )) & (~\b[5]  | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] ) | (\a[8]  ^ \a[9] )) & (~\b[6]  | (\a[10]  ^ \a[11] ) | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] )) & (~\b[4]  | (\a[9]  ^ \a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\a[8]  ^ \a[9] )));
  assign new_n78_ = \a[11]  ^ ((~new_n46_ | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] )) & (~\b[4]  | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] ) | (\a[8]  ^ \a[9] )) & (~\b[5]  | (\a[10]  ^ \a[11] ) | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] )) & (~\b[3]  | (\a[9]  ^ \a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\a[8]  ^ \a[9] )));
  assign new_n79_ = (~new_n82_ | (\a[11]  ^ (new_n81_ & (~new_n42_ | ~new_n80_)))) & ((~new_n83_ & (new_n84_ | ~new_n85_)) | (new_n82_ & (~\a[11]  ^ (new_n81_ & (~new_n42_ | ~new_n80_)))) | (~new_n82_ & (~\a[11]  | ~new_n81_ | (new_n42_ & new_n80_)) & (\a[11]  | (new_n81_ & (~new_n42_ | ~new_n80_)))));
  assign new_n80_ = (~\a[10]  | ~\a[11] ) & (\a[10]  | \a[11] ) & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] );
  assign new_n81_ = (~\b[3]  | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[4]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[2]  | (\a[9]  ^ \a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] ));
  assign new_n82_ = ((\b[0]  & (~\a[12]  | ~\a[13] ) & (\a[12]  | \a[13] ) & (\a[11]  ^ ~\a[12] )) | (\b[1]  & (~\a[13]  ^ \a[14] ) & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] )) | ((~\a[13]  | ~\a[14] ) & (\a[13]  | \a[14] ) & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ) & (\b[0]  ^ \b[1] ))) ^ (\a[14]  & \b[0]  & (\a[11]  | \a[12] ) & (~\a[11]  | ~\a[12] ));
  assign new_n83_ = \b[0]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] ) & (~\b[0]  | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[1]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\b[0]  ^ \b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\b[2]  & (\b[0]  | ~\b[1] )) | (\b[2]  & ~\b[0]  & \b[1] )) & (~\b[1]  | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[2]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[0]  | (\a[9]  ^ \a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] ));
  assign new_n84_ = \a[11]  ^ (((\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[3]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[1]  | (\a[9]  ^ \a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n85_ = (\b[0]  & (~\a[11]  | ~\a[12] ) & (\a[11]  | \a[12] )) ^ ((~\b[0]  | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[1]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\b[0]  ^ \b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\b[2]  & (\b[0]  | ~\b[1] )) | (\b[2]  & ~\b[0]  & \b[1] )) & (~\b[1]  | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[2]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & (~\b[0]  | (\a[9]  ^ \a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )));
  assign new_n86_ = ((~\b[0]  | (\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (\a[12]  ^ \a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[1]  | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[2]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\b[2]  & (\b[0]  | ~\b[1] )) | (\b[2]  & ~\b[0]  & \b[1] ))) ^ (~\a[14]  | ((~\b[0]  | (\a[12]  & \a[13] ) | (~\a[12]  & ~\a[13] ) | (~\a[11]  ^ ~\a[12] )) & (~\b[1]  | (\a[13]  ^ \a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] )) & ((\a[13]  & \a[14] ) | (~\a[13]  & ~\a[14] ) | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ) | (~\b[0]  ^ \b[1] )) & \a[14]  & (~\b[0]  | (~\a[11]  & ~\a[12] ) | (\a[11]  & \a[12] ))));
  assign new_n87_ = ~new_n72_ ^ (~new_n47_ ^ (new_n45_ ^ new_n60_));
  assign new_n88_ = \a[11]  ^ (((\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\a[8]  & \a[9] ) | (~\a[8]  & ~\a[9] ) | (~\b[8]  ^ ((\b[7]  & \b[8] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))))) & (~\b[8]  | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] ) | (\a[8]  ^ \a[9] )) & (~\b[7]  | (\a[9]  ^ \a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (\a[8]  ^ \a[9] )));
  assign new_n89_ = new_n67_ ^ ~new_n68_;
  assign new_n90_ = ~new_n91_ ^ ~\a[11] ;
  assign new_n91_ = new_n54_ ^ ((~new_n40_ & ~new_n41_) | ((new_n40_ | new_n41_) & (~new_n40_ | ~new_n41_) & ((~new_n43_ & ~new_n59_) | ((new_n43_ | new_n59_) & (~new_n43_ | ~new_n59_) & ((~new_n45_ & ~new_n60_) | (~new_n47_ & (new_n45_ | new_n60_) & (~new_n45_ | ~new_n60_)))))));
  assign new_n92_ = (new_n71_ | (~new_n73_ & new_n87_)) ^ (new_n70_ ^ ~new_n88_);
  assign new_n93_ = new_n73_ ^ ~new_n87_;
  assign new_n94_ = (~new_n96_ | new_n114_) & ((~new_n97_ & (((new_n115_ | (new_n95_ & ~new_n79_) | (~new_n95_ & new_n79_)) & (new_n99_ | (~new_n115_ & (~new_n95_ | new_n79_) & (new_n95_ | ~new_n79_)) | (new_n115_ & (~new_n95_ ^ ~new_n79_)))) | new_n97_ | new_n113_)) | (new_n96_ & ~new_n114_) | (~new_n96_ & new_n114_));
  assign new_n95_ = new_n78_ ^ ~new_n86_;
  assign new_n96_ = (new_n74_ ^ ~new_n75_) ^ ((new_n76_ & ~new_n77_) | (((~new_n78_ & new_n86_) | (~new_n79_ & (new_n78_ | ~new_n86_) & (~new_n78_ | new_n86_))) & (new_n76_ | ~new_n77_) & (~new_n76_ | new_n77_)));
  assign new_n97_ = ~new_n98_ & ((new_n76_ & ~new_n77_) | (~new_n76_ & new_n77_) | ((new_n78_ | ~new_n86_) & (new_n79_ | (~new_n78_ & new_n86_) | (new_n78_ & ~new_n86_)))) & ((new_n76_ ^ ~new_n77_) | (~new_n78_ & new_n86_) | (~new_n79_ & (new_n78_ | ~new_n86_) & (~new_n78_ | new_n86_)));
  assign new_n98_ = \a[8]  ^ (((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~\b[8]  ^ ((\b[7]  & \b[8] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))))) & (~\b[8]  | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] ) | (\a[5]  ^ \a[6] )) & (~\b[7]  | (\a[6]  ^ \a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (\a[5]  ^ \a[6] )));
  assign new_n99_ = (~new_n100_ | new_n101_) & ((new_n100_ & ~new_n101_) | (~new_n100_ & new_n101_) | ((~new_n102_ | new_n103_) & (((new_n104_ | ~new_n112_) & (new_n105_ | (~new_n104_ & new_n112_) | (new_n104_ & ~new_n112_))) | (~new_n102_ & new_n103_) | (new_n102_ & ~new_n103_))));
  assign new_n100_ = (new_n83_ | (~new_n84_ & new_n85_)) ^ (new_n82_ ^ (~\a[11]  ^ (new_n81_ & (~new_n42_ | ~new_n80_))));
  assign new_n101_ = \a[8]  ^ ((~new_n38_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] )) & (~\b[6]  | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] ) | (\a[5]  ^ \a[6] )) & (~\b[7]  | (\a[7]  ^ \a[8] ) | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] )) & (~\b[5]  | (\a[6]  ^ \a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (\a[5]  ^ \a[6] )));
  assign new_n102_ = new_n84_ ^ ~new_n85_;
  assign new_n103_ = \a[8]  ^ ((~new_n44_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] )) & (~\b[5]  | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] ) | (\a[5]  ^ \a[6] )) & (~\b[6]  | (\a[7]  ^ \a[8] ) | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] )) & (~\b[4]  | (\a[6]  ^ \a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (\a[5]  ^ \a[6] )));
  assign new_n104_ = \a[8]  ^ ((~new_n46_ | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] )) & (~\b[4]  | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] ) | (\a[5]  ^ \a[6] )) & (~\b[5]  | (\a[7]  ^ \a[8] ) | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] )) & (~\b[3]  | (\a[6]  ^ \a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (\a[5]  ^ \a[6] )));
  assign new_n105_ = (~new_n108_ | (\a[8]  ^ (new_n107_ & (~new_n42_ | ~new_n106_)))) & ((~new_n109_ & (new_n110_ | ~new_n111_)) | (new_n108_ & (~\a[8]  ^ (new_n107_ & (~new_n42_ | ~new_n106_)))) | (~new_n108_ & (~\a[8]  | ~new_n107_ | (new_n42_ & new_n106_)) & (\a[8]  | (new_n107_ & (~new_n42_ | ~new_n106_)))));
  assign new_n106_ = (~\a[7]  | ~\a[8] ) & (\a[7]  | \a[8] ) & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] );
  assign new_n107_ = (~\b[3]  | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[4]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[2]  | (\a[6]  ^ \a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] ));
  assign new_n108_ = ((\b[0]  & (~\a[9]  | ~\a[10] ) & (\a[9]  | \a[10] ) & (\a[8]  ^ ~\a[9] )) | (\b[1]  & (~\a[10]  ^ \a[11] ) & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] )) | ((~\a[10]  | ~\a[11] ) & (\a[10]  | \a[11] ) & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ) & (\b[0]  ^ \b[1] ))) ^ (\a[11]  & \b[0]  & (\a[8]  | \a[9] ) & (~\a[8]  | ~\a[9] ));
  assign new_n109_ = \b[0]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] ) & (~\b[0]  | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[1]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\b[0]  ^ \b[1] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\b[2]  & (\b[0]  | ~\b[1] )) | (\b[2]  & ~\b[0]  & \b[1] )) & (~\b[1]  | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[2]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[0]  | (\a[6]  ^ \a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] ));
  assign new_n110_ = \a[8]  ^ (((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[3]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[1]  | (\a[6]  ^ \a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n111_ = (\b[0]  & (~\a[8]  | ~\a[9] ) & (\a[8]  | \a[9] )) ^ ((~\b[0]  | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[1]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\b[0]  ^ \b[1] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\b[2]  & (\b[0]  | ~\b[1] )) | (\b[2]  & ~\b[0]  & \b[1] )) & (~\b[1]  | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[2]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & (~\b[0]  | (\a[6]  ^ \a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )));
  assign new_n112_ = (~\a[11]  | ((~\b[0]  | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[1]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\b[0]  ^ \b[1] )) & \a[11]  & (~\b[0]  | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )))) ^ ((~\b[0]  | (\a[9]  ^ \a[10] ) | (\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[1]  | (\a[9]  & \a[10] ) | (~\a[9]  & ~\a[10] ) | (~\a[8]  ^ ~\a[9] )) & (~\b[2]  | (\a[10]  ^ \a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] )) & ((\a[10]  & \a[11] ) | (~\a[10]  & ~\a[11] ) | (~\a[8]  & ~\a[9] ) | (\a[8]  & \a[9] ) | (~\b[2]  & (\b[0]  | ~\b[1] )) | (\b[2]  & ~\b[0]  & \b[1] )));
  assign new_n113_ = new_n98_ & ((~new_n76_ ^ ~new_n77_) ^ ((~new_n78_ & new_n86_) | (~new_n79_ & (new_n78_ | ~new_n86_) & (~new_n78_ | new_n86_))));
  assign new_n114_ = \a[8]  ^ (~\b[8]  | (((\a[6]  ^ \a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (\a[5]  ^ \a[6] )) & ((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | ((~\b[7]  | ~\b[8] ) & (new_n37_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))))));
  assign new_n115_ = \a[8]  ^ (((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n37_ & (~\b[7]  ^ \b[8] ))) & (~\b[7]  | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] ) | (\a[5]  ^ \a[6] )) & (~\b[8]  | (\a[7]  ^ \a[8] ) | (\a[5]  & \a[6] ) | (~\a[5]  & ~\a[6] )) & (~\b[6]  | (\a[6]  ^ \a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (\a[5]  ^ \a[6] )));
  assign new_n116_ = new_n63_ ^ (new_n39_ | new_n64_);
  assign new_n117_ = (~new_n67_ | new_n68_) & ((new_n67_ & ~new_n68_) | (~new_n67_ & new_n68_) | ((~new_n70_ | new_n88_) & ((~new_n71_ & (new_n73_ | ~new_n87_)) | (new_n70_ & ~new_n88_) | (~new_n70_ & new_n88_))));
  assign new_n118_ = ~new_n65_ ^ (\a[8]  ^ ((new_n116_ ^ \a[11] ) ^ ((new_n91_ & \a[11] ) | (~new_n117_ & (new_n91_ | \a[11] ) & (~new_n91_ | ~\a[11] )))));
  assign new_n119_ = (~new_n121_ | ~\a[5] ) & (((~\a[5]  | ((~new_n120_ | ~\a[8] ) & (new_n120_ | \a[8] ) & ((new_n92_ & \a[8] ) | ((new_n92_ | \a[8] ) & (~new_n92_ | ~\a[8] ) & ((new_n93_ & \a[8] ) | (~new_n94_ & (~new_n93_ | ~\a[8] ) & (new_n93_ | \a[8] )))))) | ((~new_n120_ ^ \a[8] ) & (~new_n92_ | ~\a[8] ) & ((~new_n92_ & ~\a[8] ) | (new_n92_ & \a[8] ) | ((~new_n93_ | ~\a[8] ) & (new_n94_ | (new_n93_ & \a[8] ) | (~new_n93_ & ~\a[8] )))))) & (((~\a[5]  | ((new_n92_ | \a[8] ) & (~new_n92_ | ~\a[8] ) & ((new_n93_ & \a[8] ) | (~new_n94_ & (~new_n93_ | ~\a[8] ) & (new_n93_ | \a[8] )))) | ((new_n92_ ^ ~\a[8] ) & (~new_n93_ | ~\a[8] ) & (new_n94_ | (new_n93_ & \a[8] ) | (~new_n93_ & ~\a[8] )))) & (new_n122_ | (\a[5]  & ((~new_n92_ & ~\a[8] ) | (new_n92_ & \a[8] ) | ((~new_n93_ | ~\a[8] ) & (new_n94_ | (new_n93_ & \a[8] ) | (~new_n93_ & ~\a[8] )))) & ((~new_n92_ ^ ~\a[8] ) | (new_n93_ & \a[8] ) | (~new_n94_ & (~new_n93_ | ~\a[8] ) & (new_n93_ | \a[8] )))) | (~\a[5]  & ((new_n92_ ^ ~\a[8] ) ^ ((new_n93_ & \a[8] ) | (~new_n94_ & (~new_n93_ | ~\a[8] ) & (new_n93_ | \a[8] ))))))) | (\a[5]  & ((new_n120_ & \a[8] ) | (~new_n120_ & ~\a[8] ) | ((~new_n92_ | ~\a[8] ) & ((~new_n92_ & ~\a[8] ) | (new_n92_ & \a[8] ) | ((~new_n93_ | ~\a[8] ) & (new_n94_ | (new_n93_ & \a[8] ) | (~new_n93_ & ~\a[8] )))))) & ((new_n120_ ^ \a[8] ) | (new_n92_ & \a[8] ) | ((new_n92_ | \a[8] ) & (~new_n92_ | ~\a[8] ) & ((new_n93_ & \a[8] ) | (~new_n94_ & (~new_n93_ | ~\a[8] ) & (new_n93_ | \a[8] )))))) | (~\a[5]  & ((~new_n120_ ^ \a[8] ) ^ ((new_n92_ & \a[8] ) | ((new_n92_ | \a[8] ) & (~new_n92_ | ~\a[8] ) & ((new_n93_ & \a[8] ) | (~new_n94_ & (~new_n93_ | ~\a[8] ) & (new_n93_ | \a[8] ))))))))) | (new_n121_ & \a[5] ) | (~new_n121_ & ~\a[5] ));
  assign new_n120_ = new_n69_ ^ ~new_n89_;
  assign new_n121_ = ((\a[8]  & (new_n69_ | ~new_n89_) & (~new_n69_ | new_n89_)) | ((~\a[8]  | (~new_n69_ & new_n89_) | (new_n69_ & ~new_n89_)) & (\a[8]  | (~new_n69_ ^ new_n89_)) & ((new_n92_ & \a[8] ) | ((~new_n92_ | ~\a[8] ) & (new_n92_ | \a[8] ) & ((new_n93_ & \a[8] ) | (~new_n94_ & (~new_n93_ | ~\a[8] ) & (new_n93_ | \a[8] ))))))) ^ (\a[8]  ^ (new_n90_ ^ (new_n66_ | (~new_n69_ & new_n89_))));
  assign new_n122_ = (~\a[5]  | (new_n94_ & ~new_n123_) | (~new_n94_ & new_n123_)) & (((~new_n124_ | ~\a[5] ) & ((~new_n124_ & ~\a[5] ) | (new_n124_ & \a[5] ) | ((~new_n126_ | ~\a[5] ) & ((~new_n126_ & ~\a[5] ) | (new_n126_ & \a[5] ) | ((~new_n127_ | ~\a[5] ) & (new_n129_ | (new_n127_ & \a[5] ) | (~new_n127_ & ~\a[5] ))))))) | (\a[5]  & (~new_n94_ | new_n123_) & (new_n94_ | ~new_n123_)) | (~\a[5]  & (~new_n94_ ^ ~new_n123_)));
  assign new_n123_ = \a[8]  ^ (new_n73_ ^ ~new_n87_);
  assign new_n124_ = new_n125_ ^ (new_n97_ | (~new_n97_ & ~new_n113_ & ((~new_n115_ & (new_n79_ | (~new_n78_ & new_n86_) | (new_n78_ & ~new_n86_)) & (~new_n79_ | (~new_n78_ ^ new_n86_))) | (~new_n99_ & (new_n115_ | (~new_n79_ & (new_n78_ | ~new_n86_) & (~new_n78_ | new_n86_)) | (new_n79_ & (new_n78_ ^ new_n86_))) & (~new_n115_ | (~new_n79_ ^ (~new_n78_ ^ new_n86_)))))));
  assign new_n125_ = ~new_n114_ ^ ((new_n74_ ^ ~new_n75_) ^ ((new_n76_ & ~new_n77_) | ((new_n76_ | ~new_n77_) & (~new_n76_ | new_n77_) & ((~new_n78_ & new_n86_) | (~new_n79_ & (new_n78_ | ~new_n86_) & (~new_n78_ | new_n86_))))));
  assign new_n126_ = (~new_n97_ & ~new_n113_) ^ ((~new_n115_ & (new_n79_ | (~new_n78_ & new_n86_) | (new_n78_ & ~new_n86_)) & (~new_n79_ | (~new_n78_ ^ new_n86_))) | (~new_n99_ & (new_n115_ | (~new_n79_ & (new_n78_ | ~new_n86_) & (~new_n78_ | new_n86_)) | (new_n79_ & (new_n78_ ^ new_n86_))) & (~new_n115_ | (~new_n79_ ^ (~new_n78_ ^ new_n86_)))));
  assign new_n127_ = new_n99_ ^ ~new_n128_;
  assign new_n128_ = ~new_n115_ ^ (~new_n79_ ^ (~new_n78_ ^ new_n86_));
  assign new_n129_ = (~new_n131_ | new_n150_) & ((new_n131_ & ~new_n150_) | (~new_n131_ & new_n150_) | (~new_n132_ & (new_n132_ | new_n134_ | ((new_n151_ | (new_n130_ & ~new_n105_) | (~new_n130_ & new_n105_)) & (new_n135_ | (~new_n151_ & (~new_n130_ | new_n105_) & (new_n130_ | ~new_n105_)) | (new_n151_ & (~new_n130_ ^ ~new_n105_)))))));
  assign new_n130_ = new_n104_ ^ ~new_n112_;
  assign new_n131_ = (new_n100_ ^ ~new_n101_) ^ ((new_n102_ & ~new_n103_) | (((~new_n104_ & new_n112_) | (~new_n105_ & (new_n104_ | ~new_n112_) & (~new_n104_ | new_n112_))) & (new_n102_ | ~new_n103_) & (~new_n102_ | new_n103_)));
  assign new_n132_ = ~new_n133_ & ((new_n102_ & ~new_n103_) | (~new_n102_ & new_n103_) | ((new_n104_ | ~new_n112_) & (new_n105_ | (~new_n104_ & new_n112_) | (new_n104_ & ~new_n112_)))) & ((new_n102_ ^ ~new_n103_) | (~new_n104_ & new_n112_) | (~new_n105_ & (new_n104_ | ~new_n112_) & (~new_n104_ | new_n112_)));
  assign new_n133_ = \a[5]  ^ (((\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~\b[8]  ^ ((\b[7]  & \b[8] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))))) & (~\b[8]  | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] ) | (\a[2]  ^ \a[3] )) & (~\b[7]  | (\a[3]  ^ \a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (\a[2]  ^ \a[3] )));
  assign new_n134_ = new_n133_ & ((~new_n102_ ^ ~new_n103_) ^ ((~new_n104_ & new_n112_) | (~new_n105_ & (new_n104_ | ~new_n112_) & (~new_n104_ | new_n112_))));
  assign new_n135_ = (~new_n136_ | new_n137_) & ((new_n136_ & ~new_n137_) | (~new_n136_ & new_n137_) | ((~new_n138_ | new_n139_) & (((new_n140_ | ~new_n149_) & (new_n143_ | (~new_n140_ & new_n149_) | (new_n140_ & ~new_n149_))) | (~new_n138_ & new_n139_) | (new_n138_ & ~new_n139_))));
  assign new_n136_ = (new_n109_ | (~new_n110_ & new_n111_)) ^ (new_n108_ ^ (~\a[8]  ^ (new_n107_ & (~new_n42_ | ~new_n106_))));
  assign new_n137_ = \a[5]  ^ ((~new_n38_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] )) & (~\b[6]  | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] ) | (\a[2]  ^ \a[3] )) & (~\b[7]  | (\a[4]  ^ \a[5] ) | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] )) & (~\b[5]  | (\a[3]  ^ \a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (\a[2]  ^ \a[3] )));
  assign new_n138_ = new_n110_ ^ ~new_n111_;
  assign new_n139_ = \a[5]  ^ ((~new_n44_ | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] )) & (~\b[5]  | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] ) | (\a[2]  ^ \a[3] )) & (~\b[6]  | (\a[4]  ^ \a[5] ) | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] )) & (~\b[4]  | (\a[3]  ^ \a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (\a[2]  ^ \a[3] )));
  assign new_n140_ = \a[5]  ^ (new_n142_ & (~new_n46_ | ~new_n141_));
  assign new_n141_ = (~\a[4]  | ~\a[5] ) & (\a[4]  | \a[5] ) & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] );
  assign new_n142_ = (~\b[4]  | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[5]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[3]  | (\a[3]  ^ \a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] ));
  assign new_n143_ = (~new_n145_ | (\a[5]  ^ (new_n144_ & (~new_n42_ | ~new_n141_)))) & ((~new_n146_ & (new_n147_ | ~new_n148_)) | (new_n145_ & (~\a[5]  ^ (new_n144_ & (~new_n42_ | ~new_n141_)))) | (~new_n145_ & (~\a[5]  | ~new_n144_ | (new_n42_ & new_n141_)) & (\a[5]  | (new_n144_ & (~new_n42_ | ~new_n141_)))));
  assign new_n144_ = (~\b[3]  | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[4]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[2]  | (\a[3]  ^ \a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] ));
  assign new_n145_ = ((\b[0]  & (~\a[6]  | ~\a[7] ) & (\a[6]  | \a[7] ) & (\a[5]  ^ ~\a[6] )) | (\b[1]  & (~\a[7]  ^ \a[8] ) & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] )) | ((~\a[7]  | ~\a[8] ) & (\a[7]  | \a[8] ) & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ) & (\b[0]  ^ \b[1] ))) ^ (\a[8]  & \b[0]  & (\a[5]  | \a[6] ) & (~\a[5]  | ~\a[6] ));
  assign new_n146_ = \b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] ) & (~\b[0]  | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[1]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\b[0]  ^ \b[1] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\b[2]  & (\b[0]  | ~\b[1] )) | (\b[2]  & ~\b[0]  & \b[1] )) & (~\b[1]  | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[2]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[0]  | (\a[3]  ^ \a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] ));
  assign new_n147_ = \a[5]  ^ (((\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[3]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[1]  | (\a[3]  ^ \a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n148_ = (\b[0]  & (~\a[5]  | ~\a[6] ) & (\a[5]  | \a[6] )) ^ ((~\b[0]  | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[1]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\b[0]  ^ \b[1] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\b[2]  & (\b[0]  | ~\b[1] )) | (\b[2]  & ~\b[0]  & \b[1] )) & (~\b[1]  | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[2]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & (~\b[0]  | (\a[3]  ^ \a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )));
  assign new_n149_ = (~\a[8]  | ((~\b[0]  | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[1]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\b[0]  ^ \b[1] )) & \a[8]  & (~\b[0]  | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )))) ^ ((~\b[0]  | (\a[6]  ^ \a[7] ) | (\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[1]  | (\a[6]  & \a[7] ) | (~\a[6]  & ~\a[7] ) | (~\a[5]  ^ ~\a[6] )) & (~\b[2]  | (\a[7]  ^ \a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] )) & ((\a[7]  & \a[8] ) | (~\a[7]  & ~\a[8] ) | (~\a[5]  & ~\a[6] ) | (\a[5]  & \a[6] ) | (~\b[2]  & (\b[0]  | ~\b[1] )) | (\b[2]  & ~\b[0]  & \b[1] )));
  assign new_n150_ = \a[5]  ^ (~\b[8]  | (((\a[3]  ^ \a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (\a[2]  ^ \a[3] )) & ((\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | ((~\b[7]  | ~\b[8] ) & (new_n37_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))))));
  assign new_n151_ = \a[5]  ^ (((\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n37_ & (~\b[7]  ^ \b[8] ))) & (~\b[7]  | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] ) | (\a[2]  ^ \a[3] )) & (~\b[8]  | (\a[4]  ^ \a[5] ) | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] )) & (~\b[6]  | (\a[3]  ^ \a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (\a[2]  ^ \a[3] )));
  assign new_n152_ = ((\a[8]  & ((new_n33_ & \a[11] ) | (~new_n33_ & ~\a[11] ) | ((~new_n116_ | ~\a[11] ) & ((~new_n116_ & ~\a[11] ) | (new_n116_ & \a[11] ) | ((~new_n91_ | ~\a[11] ) & (new_n117_ | (new_n91_ & \a[11] ) | (~new_n91_ & ~\a[11] )))))) & ((new_n33_ ^ \a[11] ) | (new_n116_ & \a[11] ) | ((new_n116_ | \a[11] ) & (~new_n116_ | ~\a[11] ) & ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] )))))) | (((\a[8]  & ((~new_n116_ & ~\a[11] ) | (new_n116_ & \a[11] ) | ((~new_n91_ | ~\a[11] ) & (new_n117_ | (new_n91_ & \a[11] ) | (~new_n91_ & ~\a[11] )))) & ((~new_n116_ ^ ~\a[11] ) | (new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] )))) | (~new_n65_ & (~\a[8]  | ((new_n116_ | \a[11] ) & (~new_n116_ | ~\a[11] ) & ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] )))) | ((new_n116_ ^ ~\a[11] ) & (~new_n91_ | ~\a[11] ) & (new_n117_ | (new_n91_ & \a[11] ) | (~new_n91_ & ~\a[11] )))) & (\a[8]  | ((~new_n116_ ^ ~\a[11] ) ^ ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] ))))))) & (~\a[8]  | ((~new_n33_ | ~\a[11] ) & (new_n33_ | \a[11] ) & ((new_n116_ & \a[11] ) | ((new_n116_ | \a[11] ) & (~new_n116_ | ~\a[11] ) & ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] )))))) | ((~new_n33_ ^ \a[11] ) & (~new_n116_ | ~\a[11] ) & ((~new_n116_ & ~\a[11] ) | (new_n116_ & \a[11] ) | ((~new_n91_ | ~\a[11] ) & (new_n117_ | (new_n91_ & \a[11] ) | (~new_n91_ & ~\a[11] )))))) & (\a[8]  | ((new_n33_ ^ \a[11] ) ^ ((new_n116_ & \a[11] ) | ((new_n116_ | \a[11] ) & (~new_n116_ | ~\a[11] ) & ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] ))))))))) ^ (\a[8]  ^ (((new_n33_ & \a[11] ) | ((~new_n33_ | ~\a[11] ) & (new_n33_ | \a[11] ) & ((new_n116_ & \a[11] ) | ((new_n116_ | \a[11] ) & (~new_n116_ | ~\a[11] ) & ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] ))))))) ^ (new_n153_ ^ \a[11] )));
  assign new_n153_ = new_n155_ ^ (new_n154_ | (new_n34_ & (new_n61_ | (new_n63_ & (new_n39_ | new_n64_)))));
  assign new_n154_ = (new_n35_ ^ \a[14] ) & ((new_n38_ & \a[16]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) | (\b[7]  & ~\a[16]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) | (\b[5]  & (~\a[14]  ^ \a[15] ) & \a[15]  & \a[16] ) | (\b[6]  & (~\a[14]  ^ \a[15] ) & (~\a[15]  | ~\a[16] ) & (\a[15]  | \a[16] )));
  assign new_n155_ = ~\a[14]  ^ ((~\b[8]  | \a[16]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] )) & (~\b[6]  | ~\a[15]  | ~\a[16]  | (\a[14]  ^ \a[15] )) & (~\b[7]  | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] ) | (\a[14]  ^ \a[15] )) & (~\a[16]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n37_ & (~\b[7]  ^ \b[8] ))));
  assign new_n156_ = (~\a[8]  | (((new_n33_ & \a[11] ) | ((~new_n33_ | ~\a[11] ) & (new_n33_ | \a[11] ) & ((new_n116_ & \a[11] ) | ((new_n116_ | \a[11] ) & (~new_n116_ | ~\a[11] ) & ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] ))))))) & (~new_n153_ | ~\a[11] ) & (new_n153_ | \a[11] )) | ((~new_n33_ | ~\a[11] ) & ((new_n33_ & \a[11] ) | (~new_n33_ & ~\a[11] ) | ((~new_n116_ | ~\a[11] ) & ((~new_n116_ & ~\a[11] ) | (new_n116_ & \a[11] ) | ((~new_n91_ | ~\a[11] ) & (new_n117_ | (new_n91_ & \a[11] ) | (~new_n91_ & ~\a[11] )))))) & (~new_n153_ ^ \a[11] ))) & (((~\a[8]  | ((~new_n33_ | ~\a[11] ) & (new_n33_ | \a[11] ) & ((new_n116_ & \a[11] ) | ((new_n116_ | \a[11] ) & (~new_n116_ | ~\a[11] ) & ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] )))))) | ((~new_n33_ ^ \a[11] ) & (~new_n116_ | ~\a[11] ) & ((~new_n116_ & ~\a[11] ) | (new_n116_ & \a[11] ) | ((~new_n91_ | ~\a[11] ) & (new_n117_ | (new_n91_ & \a[11] ) | (~new_n91_ & ~\a[11] )))))) & (((~\a[8]  | ((new_n116_ | \a[11] ) & (~new_n116_ | ~\a[11] ) & ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] )))) | ((new_n116_ ^ ~\a[11] ) & (~new_n91_ | ~\a[11] ) & (new_n117_ | (new_n91_ & \a[11] ) | (~new_n91_ & ~\a[11] )))) & (new_n65_ | (\a[8]  & ((~new_n116_ & ~\a[11] ) | (new_n116_ & \a[11] ) | ((~new_n91_ | ~\a[11] ) & (new_n117_ | (new_n91_ & \a[11] ) | (~new_n91_ & ~\a[11] )))) & ((~new_n116_ ^ ~\a[11] ) | (new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] )))) | (~\a[8]  & ((new_n116_ ^ ~\a[11] ) ^ ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] ))))))) | (\a[8]  & ((new_n33_ & \a[11] ) | (~new_n33_ & ~\a[11] ) | ((~new_n116_ | ~\a[11] ) & ((~new_n116_ & ~\a[11] ) | (new_n116_ & \a[11] ) | ((~new_n91_ | ~\a[11] ) & (new_n117_ | (new_n91_ & \a[11] ) | (~new_n91_ & ~\a[11] )))))) & ((new_n33_ ^ \a[11] ) | (new_n116_ & \a[11] ) | ((new_n116_ | \a[11] ) & (~new_n116_ | ~\a[11] ) & ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] )))))) | (~\a[8]  & ((~new_n33_ ^ \a[11] ) ^ ((new_n116_ & \a[11] ) | ((new_n116_ | \a[11] ) & (~new_n116_ | ~\a[11] ) & ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] ))))))))) | (\a[8]  & (((~new_n33_ | ~\a[11] ) & ((new_n33_ & \a[11] ) | (~new_n33_ & ~\a[11] ) | ((~new_n116_ | ~\a[11] ) & ((~new_n116_ & ~\a[11] ) | (new_n116_ & \a[11] ) | ((~new_n91_ | ~\a[11] ) & (new_n117_ | (new_n91_ & \a[11] ) | (~new_n91_ & ~\a[11] ))))))) | (new_n153_ & \a[11] ) | (~new_n153_ & ~\a[11] )) & ((new_n33_ & \a[11] ) | ((~new_n33_ | ~\a[11] ) & (new_n33_ | \a[11] ) & ((new_n116_ & \a[11] ) | ((new_n116_ | \a[11] ) & (~new_n116_ | ~\a[11] ) & ((new_n91_ & \a[11] ) | (~new_n117_ & (~new_n91_ | ~\a[11] ) & (new_n91_ | \a[11] )))))) | (new_n153_ ^ \a[11] ))) | (~\a[8]  & (((~new_n33_ | ~\a[11] ) & ((new_n33_ & \a[11] ) | (~new_n33_ & ~\a[11] ) | ((~new_n116_ | ~\a[11] ) & ((~new_n116_ & ~\a[11] ) | (new_n116_ & \a[11] ) | ((~new_n91_ | ~\a[11] ) & (new_n117_ | (new_n91_ & \a[11] ) | (~new_n91_ & ~\a[11] ))))))) ^ (new_n153_ ^ \a[11] ))));
  assign new_n157_ = (~new_n153_ | ~\a[11] ) & ((new_n153_ & \a[11] ) | (~new_n153_ & ~\a[11] ) | ((~new_n33_ | ~\a[11] ) & (((~new_n116_ | ~\a[11] ) & ((~new_n116_ & ~\a[11] ) | (new_n116_ & \a[11] ) | ((~new_n91_ | ~\a[11] ) & (new_n117_ | (new_n91_ & \a[11] ) | (~new_n91_ & ~\a[11] ))))) | (new_n33_ & \a[11] ) | (~new_n33_ & ~\a[11] ))));
  assign new_n158_ = ((\a[14]  & ((\b[8]  & ~\a[16]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) | (\b[6]  & (~\a[14]  ^ \a[15] ) & \a[15]  & \a[16] ) | (\b[7]  & (~\a[14]  ^ \a[15] ) & (~\a[15]  | ~\a[16] ) & (\a[15]  | \a[16] )) | (\a[16]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] ) & (new_n37_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )) & (~new_n37_ | (\b[7]  ^ \b[8] ))))) | (~new_n159_ & (~\a[14]  | ((~\b[8]  | \a[16]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] )) & (~\b[6]  | (\a[14]  ^ \a[15] ) | ~\a[15]  | ~\a[16] ) & (~\b[7]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\a[16]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n37_ & (~\b[7]  ^ \b[8] ))))) & (\a[14]  | (\b[8]  & ~\a[16]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) | (\b[6]  & (~\a[14]  ^ \a[15] ) & \a[15]  & \a[16] ) | (\b[7]  & (~\a[14]  ^ \a[15] ) & (~\a[15]  | ~\a[16] ) & (\a[15]  | \a[16] )) | (\a[16]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] ) & (new_n37_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )) & (~new_n37_ | (\b[7]  ^ \b[8] )))))) ^ (~\a[14]  ^ ((~\a[16]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (~\b[8]  ^ ((\b[7]  & \b[8] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))))) & (~\b[7]  | (\a[14]  ^ \a[15] ) | ~\a[15]  | ~\a[16] ) & (~\b[8]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] ))));
  assign new_n159_ = ~new_n154_ & (~new_n34_ | (~new_n61_ & (~new_n63_ | (~new_n39_ & ~new_n64_))));
  assign new_n160_ = new_n31_ ^ ~new_n161_;
  assign new_n161_ = ~new_n152_ ^ ~\a[5] ;
  assign new_n162_ = (~new_n163_ | ~\a[2] ) & (((~new_n164_ | ~\a[2] ) & ((~new_n164_ & ~\a[2] ) | (new_n164_ & \a[2] ) | ((~new_n165_ | ~\a[2] ) & (new_n168_ | (~new_n165_ & ~\a[2] ) | (new_n165_ & \a[2] ))))) | (new_n163_ & \a[2] ) | (~new_n163_ & ~\a[2] ));
  assign new_n163_ = (new_n32_ ^ \a[5] ) ^ ((new_n118_ & \a[5] ) | (~new_n119_ & (~new_n118_ | ~\a[5] ) & (new_n118_ | \a[5] )));
  assign new_n164_ = ~new_n119_ ^ (~new_n118_ ^ ~\a[5] );
  assign new_n165_ = ~new_n166_ ^ (new_n121_ ^ \a[5] );
  assign new_n166_ = (~\a[5]  | ((~new_n120_ | ~\a[8] ) & (new_n120_ | \a[8] ) & ((new_n92_ & \a[8] ) | ((~new_n92_ | ~\a[8] ) & (new_n92_ | \a[8] ) & ((new_n93_ & \a[8] ) | (~new_n94_ & new_n123_))))) | ((~new_n120_ ^ \a[8] ) & (~new_n92_ | ~\a[8] ) & ((new_n92_ & \a[8] ) | (~new_n92_ & ~\a[8] ) | ((~new_n93_ | ~\a[8] ) & (new_n94_ | ~new_n123_))))) & (((~\a[5]  | ((~new_n92_ | ~\a[8] ) & (new_n92_ | \a[8] ) & ((new_n93_ & \a[8] ) | (~new_n94_ & new_n123_))) | ((~new_n92_ ^ \a[8] ) & (~new_n93_ | ~\a[8] ) & (new_n94_ | ~new_n123_))) & (((~\a[5]  | (~new_n94_ & new_n123_) | (new_n94_ & ~new_n123_)) & (new_n167_ | (\a[5]  & (new_n94_ | ~new_n123_) & (~new_n94_ | new_n123_)) | (~\a[5]  & (new_n94_ ^ new_n123_)))) | (\a[5]  & ((new_n92_ & \a[8] ) | (~new_n92_ & ~\a[8] ) | ((~new_n93_ | ~\a[8] ) & (new_n94_ | ~new_n123_))) & ((new_n92_ ^ \a[8] ) | (new_n93_ & \a[8] ) | (~new_n94_ & new_n123_))) | (~\a[5]  & ((~new_n92_ ^ \a[8] ) ^ ((new_n93_ & \a[8] ) | (~new_n94_ & new_n123_)))))) | (\a[5]  & ((new_n120_ & \a[8] ) | (~new_n120_ & ~\a[8] ) | ((~new_n92_ | ~\a[8] ) & ((new_n92_ & \a[8] ) | (~new_n92_ & ~\a[8] ) | ((~new_n93_ | ~\a[8] ) & (new_n94_ | ~new_n123_))))) & ((new_n120_ ^ \a[8] ) | (new_n92_ & \a[8] ) | ((~new_n92_ | ~\a[8] ) & (new_n92_ | \a[8] ) & ((new_n93_ & \a[8] ) | (~new_n94_ & new_n123_))))) | (~\a[5]  & ((~new_n120_ ^ \a[8] ) ^ ((new_n92_ & \a[8] ) | ((~new_n92_ | ~\a[8] ) & (new_n92_ | \a[8] ) & ((new_n93_ & \a[8] ) | (~new_n94_ & new_n123_)))))));
  assign new_n167_ = (~new_n124_ | ~\a[5] ) & (((~new_n126_ | ~\a[5] ) & ((~new_n126_ & ~\a[5] ) | (new_n126_ & \a[5] ) | ((~new_n127_ | ~\a[5] ) & (new_n129_ | (~new_n127_ & ~\a[5] ) | (new_n127_ & \a[5] ))))) | (new_n124_ & \a[5] ) | (~new_n124_ & ~\a[5] ));
  assign new_n168_ = (~new_n169_ | ~\a[2] ) & (new_n170_ | (~new_n169_ & ~\a[2] ) | (new_n169_ & \a[2] ));
  assign new_n169_ = ((\a[5]  & ((new_n92_ & \a[8] ) | (~new_n92_ & ~\a[8] ) | ((~new_n93_ | ~\a[8] ) & (new_n94_ | ~new_n123_))) & ((new_n92_ ^ \a[8] ) | (new_n93_ & \a[8] ) | (~new_n94_ & new_n123_))) | (((\a[5]  & (new_n94_ | ~new_n123_) & (~new_n94_ | new_n123_)) | (~new_n167_ & (~\a[5]  | (~new_n94_ & new_n123_) | (new_n94_ & ~new_n123_)) & (\a[5]  | (~new_n94_ ^ new_n123_)))) & (~\a[5]  | ((~new_n92_ | ~\a[8] ) & (new_n92_ | \a[8] ) & ((new_n93_ & \a[8] ) | (~new_n94_ & new_n123_))) | ((~new_n92_ ^ \a[8] ) & (~new_n93_ | ~\a[8] ) & (new_n94_ | ~new_n123_))) & (\a[5]  | ((new_n92_ ^ \a[8] ) ^ ((new_n93_ & \a[8] ) | (~new_n94_ & new_n123_)))))) ^ (\a[5]  ^ ((new_n120_ ^ \a[8] ) ^ ((new_n92_ & \a[8] ) | ((~new_n92_ | ~\a[8] ) & (new_n92_ | \a[8] ) & ((new_n93_ & \a[8] ) | (~new_n94_ & new_n123_))))));
  assign new_n170_ = (~\a[2]  | (new_n171_ & ((\a[5]  & (new_n94_ | ~new_n123_) & (~new_n94_ | new_n123_)) | (~new_n167_ & (~\a[5]  | (~new_n94_ & new_n123_) | (new_n94_ & ~new_n123_)) & (\a[5]  | (~new_n94_ ^ new_n123_))))) | (~new_n171_ & (~\a[5]  | (~new_n94_ & new_n123_) | (new_n94_ & ~new_n123_)) & (new_n167_ | (\a[5]  & (new_n94_ | ~new_n123_) & (~new_n94_ | new_n123_)) | (~\a[5]  & (new_n94_ ^ new_n123_))))) & (((~\a[2]  | (~new_n167_ & (~\a[5]  | (~new_n94_ & new_n123_) | (new_n94_ & ~new_n123_)) & (\a[5]  | (~new_n94_ ^ new_n123_))) | (new_n167_ & (~\a[5]  ^ (~new_n94_ ^ new_n123_)))) & (((~new_n172_ | ~\a[2] ) & (new_n173_ | (~new_n172_ & ~\a[2] ) | (new_n172_ & \a[2] ))) | (\a[2]  & (new_n167_ | (\a[5]  & (new_n94_ | ~new_n123_) & (~new_n94_ | new_n123_)) | (~\a[5]  & (new_n94_ ^ new_n123_))) & (~new_n167_ | (\a[5]  ^ (~new_n94_ ^ new_n123_)))) | (~\a[2]  & (new_n167_ ^ (\a[5]  ^ (~new_n94_ ^ new_n123_)))))) | (\a[2]  & (~new_n171_ | ((~\a[5]  | (~new_n94_ & new_n123_) | (new_n94_ & ~new_n123_)) & (new_n167_ | (\a[5]  & (new_n94_ | ~new_n123_) & (~new_n94_ | new_n123_)) | (~\a[5]  & (new_n94_ ^ new_n123_))))) & (new_n171_ | (\a[5]  & (new_n94_ | ~new_n123_) & (~new_n94_ | new_n123_)) | (~new_n167_ & (~\a[5]  | (~new_n94_ & new_n123_) | (new_n94_ & ~new_n123_)) & (\a[5]  | (~new_n94_ ^ new_n123_))))) | (~\a[2]  & (~new_n171_ ^ ((\a[5]  & (new_n94_ | ~new_n123_) & (~new_n94_ | new_n123_)) | (~new_n167_ & (~\a[5]  | (~new_n94_ & new_n123_) | (new_n94_ & ~new_n123_)) & (\a[5]  | (~new_n94_ ^ new_n123_)))))));
  assign new_n171_ = \a[5]  ^ ((new_n92_ ^ \a[8] ) ^ ((new_n93_ & \a[8] ) | (~new_n94_ & (new_n93_ | \a[8] ) & (~new_n93_ | ~\a[8] ))));
  assign new_n172_ = ((new_n126_ & \a[5] ) | ((new_n126_ | \a[5] ) & (~new_n126_ | ~\a[5] ) & ((new_n127_ & \a[5] ) | (~new_n129_ & (new_n127_ | \a[5] ) & (~new_n127_ | ~\a[5] ))))) ^ (new_n124_ ^ \a[5] );
  assign new_n173_ = (~\a[2]  | ((~new_n126_ | ~\a[5] ) & (new_n126_ | \a[5] ) & ((new_n127_ & \a[5] ) | (~new_n129_ & (~new_n127_ | ~\a[5] ) & (new_n127_ | \a[5] )))) | ((~new_n126_ ^ \a[5] ) & (~new_n127_ | ~\a[5] ) & (new_n129_ | (new_n127_ & \a[5] ) | (~new_n127_ & ~\a[5] )))) & (((~\a[2]  | (~new_n129_ & (~new_n127_ | ~\a[5] ) & (new_n127_ | \a[5] )) | (new_n129_ & (~new_n127_ ^ \a[5] ))) & (((~new_n174_ | ~\a[2] ) & ((~new_n174_ & ~\a[2] ) | (new_n174_ & \a[2] ) | ((~new_n176_ | ~\a[2] ) & (new_n177_ | (new_n176_ & \a[2] ) | (~new_n176_ & ~\a[2] ))))) | (\a[2]  & (new_n129_ | (new_n127_ & \a[5] ) | (~new_n127_ & ~\a[5] )) & (~new_n129_ | (new_n127_ ^ \a[5] ))) | (~\a[2]  & (new_n129_ ^ (new_n127_ ^ \a[5] ))))) | (\a[2]  & ((new_n126_ & \a[5] ) | (~new_n126_ & ~\a[5] ) | ((~new_n127_ | ~\a[5] ) & (new_n129_ | (new_n127_ & \a[5] ) | (~new_n127_ & ~\a[5] )))) & ((new_n126_ ^ \a[5] ) | (new_n127_ & \a[5] ) | (~new_n129_ & (~new_n127_ | ~\a[5] ) & (new_n127_ | \a[5] )))) | (~\a[2]  & ((~new_n126_ ^ \a[5] ) ^ ((new_n127_ & \a[5] ) | (~new_n129_ & (~new_n127_ | ~\a[5] ) & (new_n127_ | \a[5] ))))));
  assign new_n174_ = new_n175_ ^ (new_n132_ | (~new_n132_ & ~new_n134_ & ((~new_n151_ & (new_n105_ | (~new_n104_ & new_n112_) | (new_n104_ & ~new_n112_)) & (~new_n105_ | (~new_n104_ ^ new_n112_))) | (~new_n135_ & (new_n151_ | (~new_n105_ & (new_n104_ | ~new_n112_) & (~new_n104_ | new_n112_)) | (new_n105_ & (new_n104_ ^ new_n112_))) & (~new_n151_ | (~new_n105_ ^ (~new_n104_ ^ new_n112_)))))));
  assign new_n175_ = ~new_n150_ ^ ((new_n100_ ^ ~new_n101_) ^ ((new_n102_ & ~new_n103_) | ((new_n102_ | ~new_n103_) & (~new_n102_ | new_n103_) & ((~new_n104_ & new_n112_) | (~new_n105_ & (new_n104_ | ~new_n112_) & (~new_n104_ | new_n112_))))));
  assign new_n176_ = (~new_n132_ & ~new_n134_) ^ ((~new_n151_ & (new_n105_ | (~new_n104_ & new_n112_) | (new_n104_ & ~new_n112_)) & (~new_n105_ | (~new_n104_ ^ new_n112_))) | (~new_n135_ & (new_n151_ | (~new_n105_ & (new_n104_ | ~new_n112_) & (~new_n104_ | new_n112_)) | (new_n105_ & (new_n104_ ^ new_n112_))) & (~new_n151_ | (~new_n105_ ^ (~new_n104_ ^ new_n112_)))));
  assign new_n177_ = (~\a[2]  | (new_n135_ & ~new_n178_) | (~new_n135_ & new_n178_)) & (((~new_n179_ | new_n180_) & ((~new_n179_ & new_n180_) | (new_n179_ & ~new_n180_) | (~new_n181_ & (new_n183_ | new_n181_ | new_n197_)))) | (\a[2]  & (~new_n135_ | new_n178_) & (new_n135_ | ~new_n178_)) | (~\a[2]  & (~new_n135_ ^ ~new_n178_)));
  assign new_n178_ = ~new_n151_ ^ (~new_n105_ ^ (~new_n104_ ^ new_n112_));
  assign new_n179_ = (new_n136_ ^ ~new_n137_) ^ ((new_n138_ & ~new_n139_) | (((~new_n140_ & new_n149_) | (~new_n143_ & (new_n140_ | ~new_n149_) & (~new_n140_ | new_n149_))) & (new_n138_ | ~new_n139_) & (~new_n138_ | new_n139_)));
  assign new_n180_ = \a[2]  ^ (~\b[8]  | ((new_n36_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & ((\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | \a[0]  | \a[1] )));
  assign new_n181_ = ~new_n182_ & ((new_n138_ & ~new_n139_) | (~new_n138_ & new_n139_) | ((new_n140_ | ~new_n149_) & (new_n143_ | (~new_n140_ & new_n149_) | (new_n140_ & ~new_n149_)))) & ((new_n138_ ^ ~new_n139_) | (~new_n140_ & new_n149_) | (~new_n143_ & (new_n140_ | ~new_n149_) & (~new_n140_ | new_n149_)));
  assign new_n182_ = \a[2]  ^ ((~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | (~\b[8]  ^ ((\b[7]  & \b[8] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))))) & (~\b[7]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | \a[0]  | \a[1] ) & (~\b[8]  | \a[0]  | ~\a[1] ));
  assign new_n183_ = (new_n185_ | (new_n143_ & ~new_n184_) | (~new_n143_ & new_n184_)) & (((new_n186_ | ~new_n187_) & ((~new_n186_ & new_n187_) | (new_n186_ & ~new_n187_) | ((new_n188_ | ~new_n189_) & (new_n190_ | (~new_n188_ & new_n189_) | (new_n188_ & ~new_n189_))))) | (~new_n185_ & (~new_n143_ | new_n184_) & (new_n143_ | ~new_n184_)) | (new_n185_ & (~new_n143_ ^ ~new_n184_)));
  assign new_n184_ = new_n149_ ^ (~\a[5]  ^ (new_n142_ & (~new_n46_ | ~new_n141_)));
  assign new_n185_ = \a[2]  ^ (((~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n37_ & (~\b[7]  ^ \b[8] )) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[6]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | \a[0]  | \a[1] ) & (~\b[7]  | \a[0]  | ~\a[1] ) & (~\b[8]  | ~\a[0]  | (\a[1]  ^ \a[2] )));
  assign new_n186_ = \a[2]  ^ ((~\b[5]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | \a[0]  | \a[1] ) & (~\b[6]  | \a[0]  | ~\a[1] ) & (~\b[7]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~new_n38_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )));
  assign new_n187_ = (new_n146_ | (~new_n147_ & new_n148_)) ^ (new_n145_ ^ (~\a[5]  ^ (new_n144_ & (~new_n42_ | ~new_n141_))));
  assign new_n188_ = \a[2]  ^ ((~\b[4]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | \a[0]  | \a[1] ) & (~\b[5]  | \a[0]  | ~\a[1] ) & (~\b[6]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~new_n44_ | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )));
  assign new_n189_ = new_n147_ ^ ~new_n148_;
  assign new_n190_ = (~new_n193_ | (\a[2]  ^ (new_n192_ & (~new_n46_ | ~new_n191_)))) & ((new_n193_ & (~\a[2]  ^ (new_n192_ & (~new_n46_ | ~new_n191_)))) | (~new_n193_ & (~\a[2]  | ~new_n192_ | (new_n46_ & new_n191_)) & (\a[2]  | (new_n192_ & (~new_n46_ | ~new_n191_)))) | ((new_n194_ | ~new_n195_) & (new_n196_ | (~new_n194_ & new_n195_) | (new_n194_ & ~new_n195_))));
  assign new_n191_ = \a[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] );
  assign new_n192_ = (~\b[3]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | \a[0]  | \a[1] ) & (~\b[5]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[4]  | \a[0]  | ~\a[1] );
  assign new_n193_ = (~\a[5]  | ((~\b[0]  | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[1]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\b[0]  ^ \b[1] )) & \a[5]  & (~\b[0]  | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )))) ^ ((~\b[0]  | (\a[3]  ^ \a[4] ) | (\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[1]  | (\a[3]  & \a[4] ) | (~\a[3]  & ~\a[4] ) | (~\a[2]  ^ ~\a[3] )) & (~\b[2]  | (\a[4]  ^ \a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] )) & ((\a[4]  & \a[5] ) | (~\a[4]  & ~\a[5] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  & \a[3] ) | (~\b[2]  & (\b[0]  | ~\b[1] )) | (\b[2]  & ~\b[0]  & \b[1] )));
  assign new_n194_ = \a[2]  ^ ((~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | ((~\b[3]  | ~\b[4] ) & (\b[3]  | \b[4] ) & ((\b[2]  & \b[3] ) | ((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )))) | ((~\b[3]  ^ \b[4] ) & (~\b[2]  | ~\b[3] ) & ((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )))) & (~\b[2]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | \a[0]  | \a[1] ) & (~\b[4]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[3]  | \a[0]  | ~\a[1] ));
  assign new_n195_ = ((\b[0]  & (~\a[3]  | ~\a[4] ) & (\a[3]  | \a[4] ) & (\a[2]  ^ ~\a[3] )) | (\b[1]  & (~\a[4]  ^ \a[5] ) & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] )) | ((~\a[4]  | ~\a[5] ) & (\a[4]  | \a[5] ) & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ) & (\b[0]  ^ \b[1] ))) ^ (\a[5]  & \b[0]  & (\a[2]  | \a[3] ) & (~\a[2]  | ~\a[3] ));
  assign new_n196_ = (~\b[0]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] ) | (\a[2]  ^ ((((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[3]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | \a[0]  | \a[1] ) & (~\b[2]  | \a[0]  | ~\a[1] )))) & (((~\b[0]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] )) & (~\a[2]  | (((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )) & ((\b[2]  ^ \b[3] ) | (\b[1]  & (\b[0]  | \b[2] ))) & \a[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] )) | (\b[3]  & \a[0]  & (~\a[1]  ^ \a[2] )) | (\b[1]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] ) & ~\a[0]  & ~\a[1] ) | (\b[2]  & ~\a[0]  & \a[1] )) & (\a[2]  | ((((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[3]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | \a[0]  | \a[1] ) & (~\b[2]  | \a[0]  | ~\a[1] )))) | ((\b[2]  | (~\b[0]  & \b[1] )) & (~\b[2]  | \b[0]  | ~\b[1] ) & \a[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] )) | (\b[1]  & ~\a[0]  & \a[1] ) | (\b[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] ) & ~\a[0]  & ~\a[1] ) | (\b[2]  & \a[0]  & (~\a[1]  ^ \a[2] )) | (\b[0]  & ~\a[0]  & \a[1] ) | (\b[1]  & \a[0]  & (~\a[1]  ^ \a[2] )) | ((\b[0]  ^ \b[1] ) & \a[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] )) | ~\a[2]  | (\a[0]  & \b[0] ));
  assign new_n197_ = new_n182_ & ((~new_n138_ ^ ~new_n139_) ^ ((~new_n140_ & new_n149_) | (~new_n143_ & (new_n140_ | ~new_n149_) & (~new_n140_ | new_n149_))));
  assign new_n198_ = ((~\a[5]  | (~new_n156_ & (\a[8]  | (new_n157_ ^ (~new_n158_ ^ \a[11] ))) & (~\a[8]  | (new_n157_ & (~new_n158_ ^ \a[11] )) | (~new_n157_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] )))) | (new_n156_ & (\a[8]  ^ (~new_n157_ ^ (~new_n158_ ^ \a[11] ))))) & (((~new_n152_ | ~\a[5] ) & (new_n31_ | (new_n152_ & \a[5] ) | (~new_n152_ & ~\a[5] ))) | (\a[5]  & (new_n156_ | (~\a[8]  & (~new_n157_ ^ (~new_n158_ ^ \a[11] ))) | (\a[8]  & (~new_n157_ | (new_n158_ ^ \a[11] )) & (new_n157_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] )))) & (~new_n156_ | (~\a[8]  ^ (~new_n157_ ^ (~new_n158_ ^ \a[11] ))))) | (~\a[5]  & (new_n156_ ^ (~\a[8]  ^ (~new_n157_ ^ (~new_n158_ ^ \a[11] ))))))) ^ ((\a[8]  & (~new_n157_ | (new_n158_ ^ \a[11] )) & (new_n157_ | (new_n158_ & \a[11] ) | (~new_n158_ & ~\a[11] ))) | (~new_n156_ & (\a[8]  | (new_n157_ ^ (~new_n158_ ^ \a[11] ))) & (~\a[8]  | (new_n157_ & (~new_n158_ ^ \a[11] )) | (~new_n157_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] )))));
  assign new_n199_ = ((~\a[2]  ^ (new_n31_ ^ ~new_n161_)) ^ ((new_n163_ & \a[2] ) | (((new_n164_ & \a[2] ) | ((new_n164_ | \a[2] ) & (~new_n164_ | ~\a[2] ) & ((new_n165_ & \a[2] ) | (~new_n168_ & (~new_n165_ | ~\a[2] ) & (new_n165_ | \a[2] ))))) & (~new_n163_ | ~\a[2] ) & (new_n163_ | \a[2] )))) & (((~new_n164_ | ~\a[2] ) & ((~new_n164_ & ~\a[2] ) | (new_n164_ & \a[2] ) | ((~new_n165_ | ~\a[2] ) & (new_n168_ | (new_n165_ & \a[2] ) | (~new_n165_ & ~\a[2] ))))) ^ (new_n163_ ^ \a[2] )) & ((new_n164_ ^ ~\a[2] ) ^ ((new_n165_ & \a[2] ) | (~new_n168_ & (~new_n165_ | ~\a[2] ) & (new_n165_ | \a[2] )))) & new_n200_ & (new_n168_ ^ (new_n165_ ^ \a[2] ));
  assign new_n200_ = ((~new_n169_ ^ \a[2] ) ^ ((\a[2]  & (new_n122_ | ~new_n171_) & (~new_n122_ | new_n171_)) | (((new_n201_ & \a[2] ) | ((~new_n201_ | ~\a[2] ) & (new_n201_ | \a[2] ) & ((new_n172_ & \a[2] ) | (~new_n173_ & (~new_n172_ | ~\a[2] ) & (new_n172_ | \a[2] ))))) & (~\a[2]  | (~new_n122_ & new_n171_) | (new_n122_ & ~new_n171_)) & (\a[2]  | (~new_n122_ ^ new_n171_))))) & (((~new_n201_ | ~\a[2] ) & ((new_n201_ & \a[2] ) | (~new_n201_ & ~\a[2] ) | ((~new_n172_ | ~\a[2] ) & (new_n173_ | (new_n172_ & \a[2] ) | (~new_n172_ & ~\a[2] ))))) ^ (\a[2]  ^ (~new_n122_ ^ new_n171_))) & ((new_n201_ ^ \a[2] ) | (new_n172_ & \a[2] ) | (~new_n173_ & (~new_n172_ | ~\a[2] ) & (new_n172_ | \a[2] ))) & new_n202_ & ((new_n201_ & \a[2] ) | (~new_n201_ & ~\a[2] ) | ((~new_n172_ | ~\a[2] ) & (new_n173_ | (new_n172_ & \a[2] ) | (~new_n172_ & ~\a[2] ))));
  assign new_n201_ = ~new_n167_ ^ (\a[5]  ^ (~new_n94_ ^ new_n123_));
  assign new_n202_ = (new_n206_ | (new_n203_ & \a[2] ) | ((new_n203_ | \a[2] ) & (~new_n203_ | ~\a[2] ) & ((\a[2]  & (new_n129_ | ~new_n204_) & (~new_n129_ | new_n204_)) | (~new_n205_ & (~\a[2]  | (~new_n129_ & new_n204_) | (new_n129_ & ~new_n204_)) & (\a[2]  | (~new_n129_ ^ new_n204_)))))) & (~new_n206_ | ((~new_n203_ | ~\a[2] ) & ((~new_n203_ & ~\a[2] ) | (new_n203_ & \a[2] ) | ((~\a[2]  | (~new_n129_ & new_n204_) | (new_n129_ & ~new_n204_)) & (new_n205_ | (\a[2]  & (new_n129_ | ~new_n204_) & (~new_n129_ | new_n204_)) | (~\a[2]  & (new_n129_ ^ new_n204_))))))) & ((~new_n203_ ^ ~\a[2] ) | (\a[2]  & (new_n129_ | ~new_n204_) & (~new_n129_ | new_n204_)) | (~new_n205_ & (~\a[2]  | (~new_n129_ & new_n204_) | (new_n129_ & ~new_n204_)) & (\a[2]  | (~new_n129_ ^ new_n204_)))) & ((~new_n203_ & ~\a[2] ) | (new_n203_ & \a[2] ) | ((~\a[2]  | (~new_n129_ & new_n204_) | (new_n129_ & ~new_n204_)) & (new_n205_ | (\a[2]  & (new_n129_ | ~new_n204_) & (~new_n129_ | new_n204_)) | (~\a[2]  & (new_n129_ ^ new_n204_))))) & (~new_n205_ | (\a[2]  ^ (~new_n129_ ^ new_n204_))) & new_n207_ & (new_n205_ | (\a[2]  & (new_n129_ | ~new_n204_) & (~new_n129_ | new_n204_)) | (~\a[2]  & (new_n129_ ^ new_n204_)));
  assign new_n203_ = (new_n126_ ^ \a[5] ) ^ ((~new_n129_ & new_n204_) | (new_n127_ & \a[5] ));
  assign new_n204_ = \a[5]  ^ (new_n99_ ^ ~new_n128_);
  assign new_n205_ = (~new_n174_ | ~\a[2] ) & ((new_n174_ & \a[2] ) | (~new_n174_ & ~\a[2] ) | ((~new_n176_ | ~\a[2] ) & (new_n177_ | (new_n176_ & \a[2] ) | (~new_n176_ & ~\a[2] ))));
  assign new_n206_ = \a[2]  ^ ((new_n124_ ^ \a[5] ) ^ ((new_n126_ & \a[5] ) | ((~new_n126_ | ~\a[5] ) & (new_n126_ | \a[5] ) & ((new_n127_ & \a[5] ) | (~new_n129_ & (new_n127_ | \a[5] ) & (~new_n127_ | ~\a[5] ))))));
  assign new_n207_ = ((~new_n174_ ^ \a[2] ) ^ ((new_n176_ & \a[2] ) | ((~new_n176_ | ~\a[2] ) & (new_n176_ | \a[2] ) & ((new_n208_ & \a[2] ) | ((~new_n208_ | ~\a[2] ) & (new_n208_ | \a[2] ) & ((new_n179_ & ~new_n180_) | (~new_n209_ & (new_n179_ | ~new_n180_) & (~new_n179_ | new_n180_)))))))) & ((~new_n176_ ^ \a[2] ) ^ ((new_n208_ & \a[2] ) | ((~new_n208_ | ~\a[2] ) & (new_n208_ | \a[2] ) & ((new_n179_ & ~new_n180_) | (~new_n209_ & (new_n179_ | ~new_n180_) & (~new_n179_ | new_n180_)))))) & ((new_n208_ ^ \a[2] ) | (new_n179_ & ~new_n180_) | (~new_n209_ & (new_n179_ | ~new_n180_) & (~new_n179_ | new_n180_))) & ((new_n208_ & \a[2] ) | (~new_n208_ & ~\a[2] ) | ((~new_n179_ | new_n180_) & (new_n209_ | (~new_n179_ & new_n180_) | (new_n179_ & ~new_n180_)))) & new_n210_ & (new_n209_ ^ (~new_n179_ ^ new_n180_));
  assign new_n208_ = new_n135_ ^ ~new_n178_;
  assign new_n209_ = ~new_n181_ & (new_n183_ | new_n181_ | new_n197_);
  assign new_n210_ = ((~new_n181_ & ~new_n197_) | (~new_n185_ & (new_n143_ | ~new_n184_) & (~new_n143_ | new_n184_)) | (~new_n211_ & (new_n185_ | (~new_n143_ & new_n184_) | (new_n143_ & ~new_n184_)) & (~new_n185_ | (~new_n143_ ^ new_n184_)))) & (new_n181_ | new_n197_ | ((new_n185_ | (~new_n143_ & new_n184_) | (new_n143_ & ~new_n184_)) & (new_n211_ | (~new_n185_ & (new_n143_ | ~new_n184_) & (~new_n143_ | new_n184_)) | (new_n185_ & (new_n143_ ^ new_n184_))))) & new_n212_ & (new_n211_ ^ (~new_n185_ ^ (~new_n143_ ^ new_n184_)));
  assign new_n211_ = (new_n186_ | ~new_n187_) & ((new_n186_ & ~new_n187_) | (~new_n186_ & new_n187_) | ((new_n188_ | ~new_n189_) & (new_n190_ | (~new_n188_ & new_n189_) | (new_n188_ & ~new_n189_))));
  assign new_n212_ = ((new_n186_ ^ ~new_n187_) | (~new_n188_ & new_n189_) | (~new_n190_ & (new_n188_ | ~new_n189_) & (~new_n188_ | new_n189_))) & ((new_n186_ & ~new_n187_) | (~new_n186_ & new_n187_) | ((new_n188_ | ~new_n189_) & (new_n190_ | (~new_n188_ & new_n189_) | (new_n188_ & ~new_n189_)))) & (~new_n190_ | (~new_n188_ ^ new_n189_)) & (new_n190_ | (~new_n188_ & new_n189_) | (new_n188_ & ~new_n189_)) & new_n215_ & (new_n213_ ^ new_n214_);
  assign new_n213_ = (new_n194_ | ~new_n195_) & (new_n196_ | (new_n194_ & ~new_n195_) | (~new_n194_ & new_n195_));
  assign new_n214_ = new_n193_ ^ (~\a[2]  ^ (new_n192_ & (~new_n46_ | ~new_n191_)));
  assign new_n215_ = (new_n196_ ^ (new_n194_ ^ ~new_n195_)) & ~new_n217_ & (~new_n218_ | ~new_n219_) & new_n216_ & ~new_n220_;
  assign new_n216_ = \a[0]  & \b[0] ;
  assign new_n217_ = (((\b[2]  | (~\b[0]  & \b[1] )) & (~\b[2]  | \b[0]  | ~\b[1] ) & \a[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] )) | (\b[1]  & ~\a[0]  & \a[1] ) | (\b[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] ) & ~\a[0]  & ~\a[1] ) | (\b[2]  & \a[0]  & (~\a[1]  ^ \a[2] )) | (\b[0]  & ~\a[0]  & \a[1] ) | (\b[1]  & \a[0]  & (~\a[1]  ^ \a[2] )) | ((\b[0]  ^ \b[1] ) & \a[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] )) | ~\a[2]  | (\a[0]  & \b[0] )) & (((~\b[0]  | (\a[2]  & \a[3] ) | (~\a[2]  & ~\a[3] )) & (~\a[2]  | (((\b[2]  & \b[3] ) | (~\b[2]  & ~\b[3] ) | ~\b[1]  | (~\b[0]  & ~\b[2] )) & ((\b[2]  ^ \b[3] ) | (\b[1]  & (\b[0]  | \b[2] ))) & \a[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] )) | (\b[3]  & \a[0]  & (~\a[1]  ^ \a[2] )) | (\b[1]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] ) & ~\a[0]  & ~\a[1] ) | (\b[2]  & ~\a[0]  & \a[1] )) & (\a[2]  | ((((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[3]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | \a[0]  | \a[1] ) & (~\b[2]  | \a[0]  | ~\a[1] )))) | (\b[0]  & (~\a[2]  | ~\a[3] ) & (\a[2]  | \a[3] ) & (~\a[2]  ^ ((((~\b[2]  | ~\b[3] ) & (\b[2]  | \b[3] ) & \b[1]  & (\b[0]  | \b[2] )) | ((~\b[2]  ^ \b[3] ) & (~\b[1]  | (~\b[0]  & ~\b[2] ))) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[3]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & (~\b[1]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | \a[0]  | \a[1] ) & (~\b[2]  | \a[0]  | ~\a[1] )))) | (\a[2]  & (~\a[0]  | ~\b[0]  | ((~\b[1]  | ~\a[0]  | (\a[1]  ^ \a[2] )) & ((~\b[0]  ^ \b[1] ) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ))))) | ((((~\b[2]  & (\b[0]  | ~\b[1] )) | (\b[2]  & ~\b[0]  & \b[1] ) | ~\a[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] )) & (~\b[1]  | \a[0]  | ~\a[1] ) & (~\b[0]  | (\a[1]  & \a[2] ) | (~\a[1]  & ~\a[2] ) | \a[0]  | \a[1] ) & (~\b[2]  | ~\a[0]  | (\a[1]  ^ \a[2] ))) ? ((\b[0]  & ~\a[0]  & \a[1] ) | (\b[1]  & \a[0]  & (~\a[1]  ^ \a[2] )) | ((\b[0]  ^ \b[1] ) & \a[0]  & (~\a[1]  | ~\a[2] ) & (\a[1]  | \a[2] ))) : ~\a[2] ));
  assign new_n218_ = ~\a[3]  & ~\a[4]  & ~\a[1]  & ~\a[2]  & ~\a[5]  & ~\a[8]  & ~\a[11]  & ~\a[14] ;
  assign new_n219_ = ~\a[9]  & ~\a[10]  & ~\a[6]  & ~\a[7]  & ~\a[12]  & ~\a[13]  & ~\a[15]  & ~\a[16] ;
  assign new_n220_ = ~\b[3]  & ~\b[4]  & ~\b[1]  & ~\b[2]  & ~\b[5]  & ~\b[6]  & ~\b[7]  & ~\b[8] ;
  assign new_n221_ = (\a[2]  ^ ((new_n158_ & \a[11] ) | (~new_n157_ & (~new_n158_ | ~\a[11] ) & (new_n158_ | \a[11] )))) ^ ((\a[5]  ^ \a[8] ) ^ (\a[11]  ^ \a[14] ));
  assign new_n222_ = ((~\a[14]  | ((~\a[16]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (~\b[8]  ^ ((\b[7]  & \b[8] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))))) & (~\b[7]  | (\a[14]  ^ \a[15] ) | ~\a[15]  | ~\a[16] ) & (~\b[8]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )))) & (((~\a[14]  | ((~\b[8]  | \a[16]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] )) & (~\b[6]  | (\a[14]  ^ \a[15] ) | ~\a[15]  | ~\a[16] ) & (~\b[7]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\a[16]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n37_ & (~\b[7]  ^ \b[8] ))))) & (new_n159_ | (\a[14]  & ((\b[8]  & ~\a[16]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] )) | (\b[6]  & (~\a[14]  ^ \a[15] ) & \a[15]  & \a[16] ) | (\b[7]  & (~\a[14]  ^ \a[15] ) & (~\a[15]  | ~\a[16] ) & (\a[15]  | \a[16] )) | (\a[16]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] ) & (new_n37_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] )) & (~new_n37_ | (\b[7]  ^ \b[8] ))))) | (~\a[14]  & (~\b[8]  | \a[16]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] )) & (~\b[6]  | (\a[14]  ^ \a[15] ) | ~\a[15]  | ~\a[16] ) & (~\b[7]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] )) & (~\a[16]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] )) | (new_n37_ & (~\b[7]  ^ \b[8] )))))) | (~\a[14]  & (~\a[16]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | (~\b[8]  ^ ((\b[7]  & \b[8] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))))) & (~\b[7]  | (\a[14]  ^ \a[15] ) | ~\a[15]  | ~\a[16] ) & (~\b[8]  | (\a[14]  ^ \a[15] ) | (\a[15]  & \a[16] ) | (~\a[15]  & ~\a[16] ))) | (\a[14]  & ((\a[16]  & (~\a[14]  | ~\a[15] ) & (\a[14]  | \a[15] ) & (\b[8]  ^ ((\b[7]  & \b[8] ) | (~new_n37_ & (~\b[7]  | ~\b[8] ) & (\b[7]  | \b[8] ))))) | (\b[7]  & (~\a[14]  ^ \a[15] ) & \a[15]  & \a[16] ) | (\b[8]  & (~\a[14]  ^ \a[15] ) & (~\a[15]  | ~\a[16] ) & (\a[15]  | \a[16] )))))) ^ (~\b[8]  | (((\a[14]  ^ \a[15] ) | ~\a[15]  | ~\a[16] ) & (~\a[16]  | (\a[14]  & \a[15] ) | (~\a[14]  & ~\a[15] ) | ((~\b[7]  | ~\b[8] ) & (new_n37_ | (\b[7]  & \b[8] ) | (~\b[7]  & ~\b[8] ))))));
endmodule


