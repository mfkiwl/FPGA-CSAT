// Benchmark "b14_C_sat" written by ABC on Wed Oct 26 16:38:21 2022

module b14_C_sat ( 
    DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
    DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
    DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
    DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
    DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
    DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN,
    REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN,
    REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN,
    REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN,
    REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN,
    REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN,
    REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN,
    REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN,
    IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN,
    IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN,
    IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN,
    IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN,
    IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN,
    IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN,
    IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN,
    IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN,
    IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN,
    IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN,
    IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, D_REG_1__SCAN_IN,
    D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN,
    D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
    D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
    D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
    D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
    D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
    D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
    D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
    D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
    D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
    REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
    REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
    REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
    REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
    REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
    REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
    REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
    REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
    REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
    REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
    REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
    REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
    REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
    REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
    REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
    REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
    REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
    REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
    REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
    REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
    REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
    REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
    REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
    REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
    REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
    REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
    REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
    REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
    REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
    REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
    REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
    REG2_REG_31__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_16__SCAN_IN,
    ADDR_REG_15__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_0__SCAN_IN,
    DATAO_REG_4__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_9__SCAN_IN,
    DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN,
    DATAO_REG_16__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_20__SCAN_IN,
    B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN,
    REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN,
    REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN,
    sat  );
  input  DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_,
    DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
    DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
    DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_,
    DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
    DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
    REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
    REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
    REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
    REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
    REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
    REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
    REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
    IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
    IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
    IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
    IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
    IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
    IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
    IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
    IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
    IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
    IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
    IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
    D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN,
    D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN,
    D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN,
    D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN,
    D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN,
    D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN,
    D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN,
    D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN,
    D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN,
    D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN,
    REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN,
    REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN,
    REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN,
    REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN,
    REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN,
    REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN,
    REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN,
    REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN,
    REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN,
    REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN,
    REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN,
    REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN,
    REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN,
    REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN,
    REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN,
    REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN,
    REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN,
    REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN,
    REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN,
    REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN,
    REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN,
    REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
    REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
    REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
    REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
    REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
    REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
    REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
    REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
    REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
    REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
    REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_18__SCAN_IN,
    ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_5__SCAN_IN,
    ADDR_REG_0__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_7__SCAN_IN,
    DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
    DATAO_REG_12__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_18__SCAN_IN,
    DATAO_REG_20__SCAN_IN, B_REG_SCAN_IN, REG3_REG_15__SCAN_IN,
    REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN,
    REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN;
  output sat;
  wire new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_;
  assign sat = (~new_n881_ | (~new_n241_ & new_n495_)) & ~new_n527_ & ~new_n602_ & new_n653_ & ~new_n686_ & new_n695_;
  assign new_n241_ = (~new_n248_ | ((new_n252_ & ~new_n446_) ? (~new_n242_ & ~new_n494_) : ~new_n414_)) & ~new_n362_ & (((new_n242_ | new_n494_) & new_n252_ & ~new_n446_) | new_n248_ | (new_n467_ & new_n446_));
  assign new_n242_ = new_n413_ & (~new_n387_ | (new_n412_ & (~new_n410_ | (new_n406_ & (~new_n402_ | (~new_n243_ & new_n398_))))));
  assign new_n243_ = new_n377_ & (~new_n373_ | (new_n369_ & (~new_n364_ | (new_n352_ & (~new_n386_ | (~new_n244_ & new_n383_))))));
  assign new_n244_ = new_n347_ & (~new_n343_ | (new_n338_ & (~new_n332_ | (new_n312_ & (~new_n296_ | (~new_n245_ & new_n279_))))));
  assign new_n245_ = ((((~new_n275_ ^ new_n276_) | ~new_n270_ | (~new_n275_ ^ ~new_n247_)) & (new_n272_ | ~new_n247_ | ~new_n270_) & (new_n247_ | new_n277_) & (new_n276_ | new_n270_)) | (~new_n247_ & ~new_n272_) | ~new_n270_ | (new_n247_ & ~new_n277_)) & new_n246_ & ~new_n271_ & ((~new_n275_ ^ new_n276_) | ~new_n270_ | (~new_n275_ ^ ~new_n247_) | ((new_n272_ | ~new_n247_ | ~new_n270_) & (new_n247_ | new_n277_) & (new_n276_ | new_n270_)));
  assign new_n246_ = (((new_n253_ | ~new_n247_ | ~new_n270_) & (new_n247_ | new_n261_) & (new_n260_ | new_n270_)) | (~new_n247_ & ~new_n253_) | ~new_n270_ | (new_n247_ & ~new_n261_)) & (((new_n260_ | ~new_n247_ | ~new_n270_) & (new_n267_ | new_n270_) & (new_n247_ | new_n268_)) | (~new_n247_ & ~new_n260_) | ~new_n270_ | (new_n247_ & ~new_n268_));
  assign new_n247_ = new_n248_ & new_n252_;
  assign new_n248_ = ((IR_REG_20__SCAN_IN & (~new_n251_ | ~new_n249_ | ~new_n250_)) | ~IR_REG_31__SCAN_IN | (~IR_REG_20__SCAN_IN & new_n251_ & new_n249_ & new_n250_)) & (~IR_REG_20__SCAN_IN | IR_REG_31__SCAN_IN);
  assign new_n249_ = ~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN & ~IR_REG_4__SCAN_IN & ~IR_REG_5__SCAN_IN & ~IR_REG_3__SCAN_IN & ~IR_REG_6__SCAN_IN;
  assign new_n250_ = ~IR_REG_13__SCAN_IN & ~IR_REG_11__SCAN_IN & ~IR_REG_12__SCAN_IN & ~IR_REG_7__SCAN_IN & ~IR_REG_10__SCAN_IN & ~IR_REG_8__SCAN_IN & ~IR_REG_9__SCAN_IN;
  assign new_n251_ = ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN & ~IR_REG_14__SCAN_IN & ~IR_REG_17__SCAN_IN & ~IR_REG_15__SCAN_IN & ~IR_REG_16__SCAN_IN;
  assign new_n252_ = ~IR_REG_22__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (new_n251_ & new_n249_ & new_n250_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN));
  assign new_n253_ = (~REG1_REG_4__SCAN_IN | new_n254_ | new_n257_) & (~REG0_REG_4__SCAN_IN | ~new_n254_ | new_n257_) & (~new_n259_ | new_n254_ | ~new_n257_) & (~REG2_REG_4__SCAN_IN | ~new_n254_ | ~new_n257_);
  assign new_n254_ = IR_REG_29__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_28__SCAN_IN & new_n256_ & new_n249_ & new_n250_ & new_n251_ & new_n255_));
  assign new_n255_ = ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & ~IR_REG_22__SCAN_IN & ~IR_REG_23__SCAN_IN;
  assign new_n256_ = ~IR_REG_24__SCAN_IN & ~IR_REG_25__SCAN_IN & ~IR_REG_26__SCAN_IN & ~IR_REG_27__SCAN_IN;
  assign new_n257_ = IR_REG_30__SCAN_IN ^ ((IR_REG_31__SCAN_IN & (~new_n256_ | ~new_n249_ | ~new_n250_ | ~new_n251_ | ~new_n255_)) | (~new_n258_ & IR_REG_31__SCAN_IN));
  assign new_n258_ = ~IR_REG_28__SCAN_IN & ~IR_REG_29__SCAN_IN;
  assign new_n259_ = ~REG3_REG_3__SCAN_IN ^ ~REG3_REG_4__SCAN_IN;
  assign new_n260_ = (~REG1_REG_3__SCAN_IN | new_n254_ | new_n257_) & (~REG0_REG_3__SCAN_IN | ~new_n254_ | new_n257_) & (~REG2_REG_3__SCAN_IN | ~new_n254_ | ~new_n257_) & (REG3_REG_3__SCAN_IN | new_n254_ | ~new_n257_);
  assign new_n261_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? new_n266_ : ~DATAI_4_;
  assign new_n262_ = (~IR_REG_28__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_28__SCAN_IN & new_n256_ & new_n249_ & new_n250_ & new_n251_ & new_n255_) | (IR_REG_28__SCAN_IN & (~new_n256_ | ~new_n249_ | ~new_n250_ | ~new_n251_ | ~new_n255_)));
  assign new_n263_ = IR_REG_31__SCAN_IN & (~new_n256_ | ~new_n249_ | ~new_n250_ | ~new_n251_ | ~new_n255_);
  assign new_n264_ = IR_REG_27__SCAN_IN & (IR_REG_26__SCAN_IN | IR_REG_25__SCAN_IN | IR_REG_24__SCAN_IN | ~new_n249_ | ~new_n250_ | ~new_n251_ | ~new_n255_);
  assign new_n265_ = IR_REG_27__SCAN_IN & ~IR_REG_31__SCAN_IN;
  assign new_n266_ = IR_REG_4__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_3__SCAN_IN & ~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN));
  assign new_n267_ = (~REG0_REG_2__SCAN_IN | ~new_n254_ | new_n257_) & (~REG3_REG_2__SCAN_IN | new_n254_ | ~new_n257_) & (~REG2_REG_2__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG1_REG_2__SCAN_IN | new_n254_ | new_n257_);
  assign new_n268_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? new_n269_ : ~DATAI_3_;
  assign new_n269_ = (~IR_REG_3__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_3__SCAN_IN & ~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN) | (IR_REG_3__SCAN_IN & (IR_REG_2__SCAN_IN | IR_REG_0__SCAN_IN | IR_REG_1__SCAN_IN)));
  assign new_n270_ = IR_REG_23__SCAN_IN ^ ((IR_REG_31__SCAN_IN & (~new_n251_ | ~new_n249_ | ~new_n250_ | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN)) | (IR_REG_22__SCAN_IN & IR_REG_31__SCAN_IN));
  assign new_n271_ = ((~new_n267_ & new_n247_ & new_n270_) | (~new_n272_ & ~new_n270_) | (~new_n247_ & new_n273_)) & (new_n247_ | new_n267_) & new_n270_ & (~new_n247_ | ~new_n273_);
  assign new_n272_ = (~REG1_REG_1__SCAN_IN | new_n254_ | new_n257_) & (~REG2_REG_1__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG0_REG_1__SCAN_IN | ~new_n254_ | new_n257_) & (~REG3_REG_1__SCAN_IN | new_n254_ | ~new_n257_);
  assign new_n273_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? new_n274_ : DATAI_2_;
  assign new_n274_ = IR_REG_31__SCAN_IN ? (~IR_REG_2__SCAN_IN ^ (~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN)) : IR_REG_2__SCAN_IN;
  assign new_n275_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? ~IR_REG_0__SCAN_IN : ~DATAI_0_;
  assign new_n276_ = (~REG1_REG_0__SCAN_IN | new_n254_ | new_n257_) & (~REG0_REG_0__SCAN_IN | ~new_n254_ | new_n257_) & (~REG3_REG_0__SCAN_IN | new_n254_ | ~new_n257_) & (~REG2_REG_0__SCAN_IN | ~new_n254_ | ~new_n257_);
  assign new_n277_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? ~new_n278_ : ~DATAI_1_;
  assign new_n278_ = ~IR_REG_1__SCAN_IN ^ (~IR_REG_0__SCAN_IN | ~IR_REG_31__SCAN_IN);
  assign new_n279_ = (~new_n246_ | ~new_n280_) & ~new_n281_ & new_n282_ & new_n286_;
  assign new_n280_ = (new_n267_ | ~new_n247_ | ~new_n270_) & (new_n272_ | new_n270_) & (new_n247_ | ~new_n273_) & ((~new_n247_ & ~new_n267_) | ~new_n270_ | (new_n247_ & new_n273_));
  assign new_n281_ = (((new_n253_ | ~new_n247_ | ~new_n270_) & (new_n247_ | new_n261_) & (new_n260_ | new_n270_)) | (~new_n247_ & ~new_n253_) | ~new_n270_ | (new_n247_ & ~new_n261_)) & (new_n260_ | ~new_n247_ | ~new_n270_) & (new_n267_ | new_n270_) & (new_n247_ | new_n268_) & ((~new_n247_ & ~new_n260_) | ~new_n270_ | (new_n247_ & ~new_n268_));
  assign new_n282_ = ((~new_n253_ & new_n247_ & new_n270_) | (~new_n247_ & ~new_n261_) | (~new_n260_ & ~new_n270_) | ((new_n247_ | new_n253_) & new_n270_ & (~new_n247_ | new_n261_))) & ((~new_n283_ & new_n247_ & new_n270_) | (~new_n247_ & ~new_n284_) | (~new_n253_ & ~new_n270_) | (new_n270_ & (~new_n247_ | new_n284_) & (new_n247_ | new_n283_)));
  assign new_n283_ = (~REG1_REG_5__SCAN_IN | new_n254_ | new_n257_) & (~REG2_REG_5__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG0_REG_5__SCAN_IN | ~new_n254_ | new_n257_) & (new_n254_ | ~new_n257_ | (REG3_REG_5__SCAN_IN & REG3_REG_3__SCAN_IN & REG3_REG_4__SCAN_IN) | (~REG3_REG_5__SCAN_IN & (~REG3_REG_3__SCAN_IN | ~REG3_REG_4__SCAN_IN)));
  assign new_n284_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? ~new_n285_ : ~DATAI_5_;
  assign new_n285_ = IR_REG_5__SCAN_IN ^ ((IR_REG_31__SCAN_IN & (IR_REG_3__SCAN_IN | IR_REG_2__SCAN_IN | IR_REG_0__SCAN_IN | IR_REG_1__SCAN_IN)) | (IR_REG_4__SCAN_IN & IR_REG_31__SCAN_IN));
  assign new_n286_ = ((~new_n247_ & ~new_n287_) | (~new_n289_ & ~new_n270_) | (~new_n291_ & new_n247_ & new_n270_) | ((~new_n247_ | new_n287_) & new_n270_ & (new_n247_ | new_n291_))) & ((~new_n289_ & new_n247_ & new_n270_) | (~new_n283_ & ~new_n270_) | (~new_n247_ & new_n293_) | ((new_n247_ | new_n289_) & new_n270_ & (~new_n247_ | ~new_n293_)));
  assign new_n287_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? ~new_n288_ : ~DATAI_7_;
  assign new_n288_ = ~IR_REG_7__SCAN_IN ^ (new_n249_ | ~IR_REG_31__SCAN_IN);
  assign new_n289_ = (~REG1_REG_6__SCAN_IN | new_n254_ | new_n257_) & (~REG0_REG_6__SCAN_IN | ~new_n254_ | new_n257_) & (~new_n290_ | new_n254_ | ~new_n257_) & (~REG2_REG_6__SCAN_IN | ~new_n254_ | ~new_n257_);
  assign new_n290_ = REG3_REG_6__SCAN_IN ^ (REG3_REG_5__SCAN_IN & REG3_REG_3__SCAN_IN & REG3_REG_4__SCAN_IN);
  assign new_n291_ = (~REG2_REG_7__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG1_REG_7__SCAN_IN | new_n254_ | new_n257_) & (~REG0_REG_7__SCAN_IN | ~new_n254_ | new_n257_) & (new_n254_ | ~new_n257_ | (new_n292_ & REG3_REG_7__SCAN_IN) | (~new_n292_ & ~REG3_REG_7__SCAN_IN));
  assign new_n292_ = REG3_REG_6__SCAN_IN & REG3_REG_5__SCAN_IN & REG3_REG_3__SCAN_IN & REG3_REG_4__SCAN_IN;
  assign new_n293_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? new_n294_ : DATAI_6_;
  assign new_n294_ = IR_REG_31__SCAN_IN ? (~new_n249_ & ~new_n295_) : IR_REG_6__SCAN_IN;
  assign new_n295_ = IR_REG_6__SCAN_IN & (IR_REG_4__SCAN_IN | IR_REG_5__SCAN_IN | IR_REG_3__SCAN_IN | IR_REG_2__SCAN_IN | IR_REG_0__SCAN_IN | IR_REG_1__SCAN_IN);
  assign new_n296_ = (new_n297_ | ((new_n247_ | new_n287_) & (new_n289_ | new_n270_) & (new_n291_ | ~new_n247_ | ~new_n270_) & ((new_n247_ & ~new_n287_) | ~new_n270_ | (~new_n247_ & ~new_n291_)))) & new_n298_ & ~new_n309_ & (((new_n247_ | new_n287_) & (new_n289_ | new_n270_) & (new_n291_ | ~new_n247_ | ~new_n270_)) | (new_n247_ & ~new_n287_) | ~new_n270_ | (~new_n247_ & ~new_n291_));
  assign new_n297_ = (((new_n289_ | ~new_n247_ | ~new_n270_) & (new_n283_ | new_n270_) & (new_n247_ | ~new_n293_)) | (~new_n247_ & ~new_n289_) | ~new_n270_ | (new_n247_ & new_n293_)) & (((new_n289_ | ~new_n247_ | ~new_n270_) & (new_n283_ | new_n270_) & (new_n247_ | ~new_n293_) & ((~new_n247_ & ~new_n289_) | ~new_n270_ | (new_n247_ & new_n293_))) | ((new_n283_ | ~new_n247_ | ~new_n270_) & (new_n247_ | new_n284_) & (new_n253_ | new_n270_)) | ~new_n270_ | (new_n247_ & ~new_n284_) | (~new_n247_ & ~new_n283_));
  assign new_n298_ = (((new_n299_ | ~new_n247_ | ~new_n270_) & (new_n247_ | new_n303_) & (new_n301_ | new_n270_)) | (~new_n247_ & ~new_n299_) | ~new_n270_ | (new_n247_ & ~new_n303_)) & (((new_n301_ | ~new_n247_ | ~new_n270_) & (new_n306_ | new_n270_) & (new_n247_ | new_n307_)) | (~new_n247_ & ~new_n301_) | ~new_n270_ | (new_n247_ & ~new_n307_));
  assign new_n299_ = (~REG1_REG_10__SCAN_IN | new_n254_ | new_n257_) & (new_n254_ | ~new_n257_ | (new_n300_ & REG3_REG_10__SCAN_IN) | (~new_n300_ & ~REG3_REG_10__SCAN_IN)) & (~REG2_REG_10__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG0_REG_10__SCAN_IN | ~new_n254_ | new_n257_);
  assign new_n300_ = REG3_REG_9__SCAN_IN & REG3_REG_8__SCAN_IN & REG3_REG_7__SCAN_IN & REG3_REG_6__SCAN_IN & REG3_REG_5__SCAN_IN & REG3_REG_3__SCAN_IN & REG3_REG_4__SCAN_IN;
  assign new_n301_ = (~REG1_REG_9__SCAN_IN | new_n254_ | new_n257_) & (new_n254_ | ~new_n257_ | (new_n302_ & REG3_REG_9__SCAN_IN) | (~new_n302_ & ~REG3_REG_9__SCAN_IN)) & (~REG2_REG_9__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG0_REG_9__SCAN_IN | ~new_n254_ | new_n257_);
  assign new_n302_ = REG3_REG_8__SCAN_IN & new_n292_ & REG3_REG_7__SCAN_IN;
  assign new_n303_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? new_n304_ : ~DATAI_10_;
  assign new_n304_ = IR_REG_10__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (new_n305_ & new_n249_ & ~IR_REG_7__SCAN_IN));
  assign new_n305_ = ~IR_REG_8__SCAN_IN & ~IR_REG_9__SCAN_IN;
  assign new_n306_ = (~REG1_REG_8__SCAN_IN | new_n254_ | new_n257_) & (~REG2_REG_8__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG0_REG_8__SCAN_IN | ~new_n254_ | new_n257_) & (new_n254_ | ~new_n257_ | (REG3_REG_8__SCAN_IN & new_n292_ & REG3_REG_7__SCAN_IN) | (~REG3_REG_8__SCAN_IN & (~new_n292_ | ~REG3_REG_7__SCAN_IN)));
  assign new_n307_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? new_n308_ : ~DATAI_9_;
  assign new_n308_ = (~IR_REG_9__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (new_n249_ & ~IR_REG_7__SCAN_IN & ~IR_REG_8__SCAN_IN & ~IR_REG_9__SCAN_IN) | (IR_REG_9__SCAN_IN & (IR_REG_8__SCAN_IN | ~new_n249_ | IR_REG_7__SCAN_IN)));
  assign new_n309_ = ((~new_n306_ & new_n247_ & new_n270_) | (~new_n291_ & ~new_n270_) | (~new_n247_ & new_n310_)) & (new_n247_ | new_n306_) & new_n270_ & (~new_n247_ | ~new_n310_);
  assign new_n310_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? new_n311_ : DATAI_8_;
  assign new_n311_ = IR_REG_31__SCAN_IN ? (~IR_REG_8__SCAN_IN ^ (new_n249_ & ~IR_REG_7__SCAN_IN)) : IR_REG_8__SCAN_IN;
  assign new_n312_ = (~new_n316_ | new_n313_ | (~new_n314_ & new_n315_)) & ~new_n317_ & ~new_n324_ & (new_n313_ | ~new_n314_ | new_n315_) & ~new_n328_ & ~new_n331_;
  assign new_n313_ = ((~new_n299_ & new_n247_ & new_n270_) | (~new_n247_ & ~new_n303_) | (~new_n301_ & ~new_n270_)) & (new_n247_ | new_n299_) & new_n270_ & (~new_n247_ | new_n303_);
  assign new_n314_ = (new_n301_ | ~new_n247_ | ~new_n270_) & (new_n247_ | new_n307_) & (new_n306_ | new_n270_);
  assign new_n315_ = (new_n247_ | new_n301_) & new_n270_ & (~new_n247_ | new_n307_);
  assign new_n316_ = (new_n306_ | ~new_n247_ | ~new_n270_) & (new_n291_ | new_n270_) & (new_n247_ | ~new_n310_) & ((~new_n247_ & ~new_n306_) | ~new_n270_ | (new_n247_ & new_n310_));
  assign new_n317_ = (new_n247_ | new_n318_) & (new_n320_ | new_n270_) & (new_n322_ | ~new_n247_ | ~new_n270_) & ((~new_n247_ & ~new_n322_) | ~new_n270_ | (new_n247_ & ~new_n318_));
  assign new_n318_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? new_n319_ : ~DATAI_13_;
  assign new_n319_ = (~IR_REG_13__SCAN_IN | IR_REG_31__SCAN_IN) & ((IR_REG_13__SCAN_IN & (IR_REG_12__SCAN_IN | IR_REG_11__SCAN_IN | IR_REG_10__SCAN_IN | ~new_n305_ | ~new_n249_ | IR_REG_7__SCAN_IN)) | ~IR_REG_31__SCAN_IN | (new_n249_ & ~IR_REG_13__SCAN_IN & ~IR_REG_11__SCAN_IN & ~IR_REG_12__SCAN_IN & new_n305_ & ~IR_REG_7__SCAN_IN & ~IR_REG_10__SCAN_IN));
  assign new_n320_ = (~REG2_REG_12__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG1_REG_12__SCAN_IN | new_n254_ | new_n257_) & (~REG0_REG_12__SCAN_IN | ~new_n254_ | new_n257_) & (new_n254_ | ~new_n257_ | (REG3_REG_12__SCAN_IN & new_n321_ & REG3_REG_11__SCAN_IN) | (~REG3_REG_12__SCAN_IN & (~new_n321_ | ~REG3_REG_11__SCAN_IN)));
  assign new_n321_ = REG3_REG_10__SCAN_IN & REG3_REG_9__SCAN_IN & REG3_REG_8__SCAN_IN & REG3_REG_7__SCAN_IN & REG3_REG_6__SCAN_IN & REG3_REG_5__SCAN_IN & REG3_REG_3__SCAN_IN & REG3_REG_4__SCAN_IN;
  assign new_n322_ = (~REG1_REG_13__SCAN_IN | new_n254_ | new_n257_) & (new_n254_ | ~new_n257_ | (new_n323_ & REG3_REG_13__SCAN_IN) | (~new_n323_ & ~REG3_REG_13__SCAN_IN)) & (~REG2_REG_13__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG0_REG_13__SCAN_IN | ~new_n254_ | new_n257_);
  assign new_n323_ = REG3_REG_12__SCAN_IN & new_n321_ & REG3_REG_11__SCAN_IN;
  assign new_n324_ = (new_n247_ | ~new_n325_) & (new_n327_ | new_n270_) & (new_n320_ | ~new_n247_ | ~new_n270_) & ((~new_n247_ & ~new_n320_) | ~new_n270_ | (new_n247_ & new_n325_));
  assign new_n325_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? new_n326_ : DATAI_12_;
  assign new_n326_ = IR_REG_31__SCAN_IN ? (~IR_REG_12__SCAN_IN ^ (~IR_REG_11__SCAN_IN & ~IR_REG_10__SCAN_IN & new_n305_ & new_n249_ & ~IR_REG_7__SCAN_IN)) : IR_REG_12__SCAN_IN;
  assign new_n327_ = (~REG1_REG_11__SCAN_IN | new_n254_ | new_n257_) & (~REG2_REG_11__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG0_REG_11__SCAN_IN | ~new_n254_ | new_n257_) & (new_n254_ | ~new_n257_ | (new_n321_ & REG3_REG_11__SCAN_IN) | (~new_n321_ & ~REG3_REG_11__SCAN_IN));
  assign new_n328_ = (new_n327_ | ~new_n247_ | ~new_n270_) & (new_n247_ | new_n329_) & (new_n299_ | new_n270_) & ((~new_n247_ & ~new_n327_) | ~new_n270_ | (new_n247_ & ~new_n329_));
  assign new_n329_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? ~new_n330_ : ~DATAI_11_;
  assign new_n330_ = ~IR_REG_11__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_10__SCAN_IN & new_n305_ & new_n249_ & ~IR_REG_7__SCAN_IN));
  assign new_n331_ = (new_n299_ | ~new_n247_ | ~new_n270_) & (new_n247_ | new_n303_) & (new_n301_ | new_n270_) & ((~new_n247_ & ~new_n299_) | ~new_n270_ | (new_n247_ & ~new_n303_));
  assign new_n332_ = (~new_n333_ | new_n317_ | ((new_n247_ | ~new_n325_) & (new_n327_ | new_n270_) & (new_n320_ | ~new_n247_ | ~new_n270_) & ((~new_n247_ & ~new_n320_) | ~new_n270_ | (new_n247_ & new_n325_)))) & new_n334_ & (new_n317_ | ((new_n247_ | ~new_n325_) & (new_n327_ | new_n270_) & (new_n320_ | ~new_n247_ | ~new_n270_)) | (~new_n247_ & ~new_n320_) | ~new_n270_ | (new_n247_ & new_n325_));
  assign new_n333_ = ((~new_n327_ & new_n247_ & new_n270_) | (~new_n247_ & ~new_n329_) | (~new_n299_ & ~new_n270_)) & (new_n247_ | new_n327_) & new_n270_ & (~new_n247_ | new_n329_);
  assign new_n334_ = (~new_n270_ | (new_n247_ & ~new_n336_) | (~new_n247_ & ~new_n335_) | ((new_n335_ | ~new_n247_ | ~new_n270_) & (new_n247_ | new_n336_) & (new_n322_ | new_n270_))) & (((new_n247_ | new_n318_) & (new_n320_ | new_n270_) & (new_n322_ | ~new_n247_ | ~new_n270_)) | (~new_n247_ & ~new_n322_) | ~new_n270_ | (new_n247_ & ~new_n318_));
  assign new_n335_ = ((~REG3_REG_14__SCAN_IN & (~new_n323_ | ~REG3_REG_13__SCAN_IN)) | new_n254_ | ~new_n257_ | (REG3_REG_14__SCAN_IN & new_n323_ & REG3_REG_13__SCAN_IN)) & (~REG1_REG_14__SCAN_IN | new_n254_ | new_n257_) & (~REG2_REG_14__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG0_REG_14__SCAN_IN | ~new_n254_ | new_n257_);
  assign new_n336_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? new_n337_ : ~DATAI_14_;
  assign new_n337_ = IR_REG_14__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (new_n249_ & new_n250_));
  assign new_n338_ = ((~new_n335_ & new_n247_ & new_n270_) | (~new_n247_ & ~new_n336_) | (~new_n322_ & ~new_n270_) | (new_n270_ & (~new_n247_ | new_n336_) & (new_n247_ | new_n335_))) & ((new_n270_ & (~new_n247_ | new_n341_) & (new_n247_ | new_n339_)) | (~new_n335_ & ~new_n270_) | (~new_n247_ & ~new_n341_) | (~new_n339_ & new_n247_ & new_n270_));
  assign new_n339_ = (new_n254_ | ~new_n257_ | (new_n340_ & REG3_REG_15__SCAN_IN) | (~new_n340_ & ~REG3_REG_15__SCAN_IN)) & (~REG0_REG_15__SCAN_IN | ~new_n254_ | new_n257_) & (~REG1_REG_15__SCAN_IN | new_n254_ | new_n257_) & (~REG2_REG_15__SCAN_IN | ~new_n254_ | ~new_n257_);
  assign new_n340_ = REG3_REG_14__SCAN_IN & REG3_REG_13__SCAN_IN & REG3_REG_12__SCAN_IN & new_n321_ & REG3_REG_11__SCAN_IN;
  assign new_n341_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? ~new_n342_ : ~DATAI_15_;
  assign new_n342_ = IR_REG_31__SCAN_IN ? (~IR_REG_15__SCAN_IN ^ (~IR_REG_14__SCAN_IN & new_n249_ & new_n250_)) : IR_REG_15__SCAN_IN;
  assign new_n343_ = (~new_n270_ | (new_n247_ & ~new_n341_) | (~new_n247_ & ~new_n339_) | ((new_n335_ | new_n270_) & (new_n247_ | new_n341_) & (new_n339_ | ~new_n247_ | ~new_n270_))) & (~new_n270_ | (new_n247_ & ~new_n345_) | (~new_n247_ & ~new_n344_) | ((new_n344_ | ~new_n247_ | ~new_n270_) & (new_n339_ | new_n270_) & (new_n247_ | new_n345_)));
  assign new_n344_ = ((~REG3_REG_16__SCAN_IN & (~new_n340_ | ~REG3_REG_15__SCAN_IN)) | new_n254_ | ~new_n257_ | (REG3_REG_16__SCAN_IN & new_n340_ & REG3_REG_15__SCAN_IN)) & (~REG2_REG_16__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG1_REG_16__SCAN_IN | new_n254_ | new_n257_) & (~REG0_REG_16__SCAN_IN | ~new_n254_ | new_n257_);
  assign new_n345_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? ~new_n346_ : ~DATAI_16_;
  assign new_n346_ = IR_REG_31__SCAN_IN ? ((~IR_REG_16__SCAN_IN | (~IR_REG_15__SCAN_IN & ~IR_REG_14__SCAN_IN & new_n249_ & new_n250_)) & (IR_REG_15__SCAN_IN | IR_REG_16__SCAN_IN | IR_REG_14__SCAN_IN | ~new_n249_ | ~new_n250_)) : IR_REG_16__SCAN_IN;
  assign new_n347_ = ((~new_n344_ & new_n247_ & new_n270_) | (~new_n247_ & ~new_n345_) | (~new_n339_ & ~new_n270_) | (new_n270_ & (~new_n247_ | new_n345_) & (new_n247_ | new_n344_))) & ((new_n270_ & (~new_n247_ | new_n350_) & (new_n247_ | new_n348_)) | (~new_n348_ & new_n247_ & new_n270_) | (~new_n344_ & ~new_n270_) | (~new_n247_ & ~new_n350_));
  assign new_n348_ = (new_n254_ | ~new_n257_ | (new_n349_ & REG3_REG_17__SCAN_IN) | (~new_n349_ & ~REG3_REG_17__SCAN_IN)) & (~REG2_REG_17__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG1_REG_17__SCAN_IN | new_n254_ | new_n257_) & (~REG0_REG_17__SCAN_IN | ~new_n254_ | new_n257_);
  assign new_n349_ = REG3_REG_16__SCAN_IN & REG3_REG_15__SCAN_IN & REG3_REG_14__SCAN_IN & REG3_REG_13__SCAN_IN & REG3_REG_12__SCAN_IN & new_n321_ & REG3_REG_11__SCAN_IN;
  assign new_n350_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? new_n351_ : ~DATAI_17_;
  assign new_n351_ = (~IR_REG_17__SCAN_IN | IR_REG_31__SCAN_IN) & ((IR_REG_17__SCAN_IN & (IR_REG_15__SCAN_IN | IR_REG_16__SCAN_IN | IR_REG_14__SCAN_IN | ~new_n249_ | ~new_n250_)) | ~IR_REG_31__SCAN_IN | (new_n249_ & new_n250_ & ~IR_REG_15__SCAN_IN & ~IR_REG_16__SCAN_IN & ~IR_REG_14__SCAN_IN & ~IR_REG_17__SCAN_IN));
  assign new_n352_ = (((new_n360_ | ~new_n247_ | ~new_n270_) & (new_n359_ | new_n270_) & (new_n247_ | new_n361_)) | (~new_n247_ & ~new_n360_) | ~new_n270_ | (new_n247_ & ~new_n361_)) & (((new_n353_ | ~new_n247_ | ~new_n270_) & (new_n360_ | new_n270_) & (~new_n357_ | new_n247_)) | (~new_n353_ & ~new_n247_) | ~new_n270_ | (new_n357_ & new_n247_));
  assign new_n353_ = ~new_n354_ & new_n356_;
  assign new_n354_ = (REG3_REG_20__SCAN_IN | (REG3_REG_19__SCAN_IN & new_n355_ & REG3_REG_18__SCAN_IN)) & ~new_n254_ & new_n257_ & (~REG3_REG_20__SCAN_IN | ~REG3_REG_19__SCAN_IN | ~new_n355_ | ~REG3_REG_18__SCAN_IN);
  assign new_n355_ = REG3_REG_17__SCAN_IN & REG3_REG_16__SCAN_IN & REG3_REG_15__SCAN_IN & REG3_REG_14__SCAN_IN & REG3_REG_13__SCAN_IN & REG3_REG_12__SCAN_IN & new_n321_ & REG3_REG_11__SCAN_IN;
  assign new_n356_ = (~REG0_REG_20__SCAN_IN | ~new_n254_ | new_n257_) & (~REG2_REG_20__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG1_REG_20__SCAN_IN | new_n254_ | new_n257_);
  assign new_n357_ = ~new_n358_ & DATAI_20_;
  assign new_n358_ = new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_);
  assign new_n359_ = (new_n254_ | ~new_n257_ | (new_n355_ & REG3_REG_18__SCAN_IN) | (~new_n355_ & ~REG3_REG_18__SCAN_IN)) & (~REG0_REG_18__SCAN_IN | ~new_n254_ | new_n257_) & (~REG1_REG_18__SCAN_IN | new_n254_ | new_n257_) & (~REG2_REG_18__SCAN_IN | ~new_n254_ | ~new_n257_);
  assign new_n360_ = ((~REG3_REG_19__SCAN_IN & (~new_n355_ | ~REG3_REG_18__SCAN_IN)) | new_n254_ | ~new_n257_ | (REG3_REG_19__SCAN_IN & new_n355_ & REG3_REG_18__SCAN_IN)) & (~REG1_REG_19__SCAN_IN | new_n254_ | new_n257_) & (~REG2_REG_19__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG0_REG_19__SCAN_IN | ~new_n254_ | new_n257_);
  assign new_n361_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? ~new_n362_ : ~DATAI_19_;
  assign new_n362_ = (~IR_REG_19__SCAN_IN | ~IR_REG_31__SCAN_IN | (~IR_REG_18__SCAN_IN & new_n363_ & new_n249_ & new_n250_)) & (IR_REG_19__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | ~new_n249_ | ~new_n250_ | ~new_n363_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN);
  assign new_n363_ = ~IR_REG_14__SCAN_IN & ~IR_REG_17__SCAN_IN & ~IR_REG_15__SCAN_IN & ~IR_REG_16__SCAN_IN;
  assign new_n364_ = ((~new_n353_ & new_n247_ & new_n270_) | (~new_n360_ & ~new_n270_) | (new_n357_ & ~new_n247_) | ((new_n353_ | new_n247_) & new_n270_ & (~new_n357_ | ~new_n247_))) & ((~new_n365_ & new_n247_ & new_n270_) | (~new_n247_ & new_n368_) | (~new_n353_ & ~new_n270_) | ((new_n365_ | new_n247_) & new_n270_ & (~new_n247_ | ~new_n368_)));
  assign new_n365_ = new_n367_ & ((~REG3_REG_21__SCAN_IN & (~REG3_REG_20__SCAN_IN | ~REG3_REG_19__SCAN_IN | ~new_n355_ | ~REG3_REG_18__SCAN_IN)) | ~new_n366_ | (REG3_REG_21__SCAN_IN & REG3_REG_20__SCAN_IN & REG3_REG_19__SCAN_IN & new_n355_ & REG3_REG_18__SCAN_IN));
  assign new_n366_ = ~new_n254_ & new_n257_;
  assign new_n367_ = (~REG0_REG_21__SCAN_IN | ~new_n254_ | new_n257_) & (~REG2_REG_21__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG1_REG_21__SCAN_IN | new_n254_ | new_n257_);
  assign new_n368_ = DATAI_21_ & (~new_n262_ | new_n265_ | (new_n263_ & ~new_n264_));
  assign new_n369_ = (((new_n365_ | ~new_n247_ | ~new_n270_) & (new_n353_ | new_n270_) & (new_n247_ | new_n358_ | ~DATAI_21_)) | (~new_n365_ & ~new_n247_) | ~new_n270_ | (new_n247_ & ~new_n358_ & DATAI_21_)) & (((new_n370_ | ~new_n247_ | ~new_n270_) & (new_n247_ | new_n358_ | ~DATAI_22_) & (new_n365_ | new_n270_)) | (~new_n370_ & ~new_n247_) | ~new_n270_ | (new_n247_ & ~new_n358_ & DATAI_22_));
  assign new_n370_ = new_n372_ & ((~new_n371_ & ~REG3_REG_22__SCAN_IN) | ~new_n366_ | (new_n371_ & REG3_REG_22__SCAN_IN));
  assign new_n371_ = REG3_REG_21__SCAN_IN & REG3_REG_20__SCAN_IN & REG3_REG_19__SCAN_IN & new_n355_ & REG3_REG_18__SCAN_IN;
  assign new_n372_ = (~REG0_REG_22__SCAN_IN | ~new_n254_ | new_n257_) & (~REG2_REG_22__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG1_REG_22__SCAN_IN | new_n254_ | new_n257_);
  assign new_n373_ = ((~new_n370_ & new_n247_ & new_n270_) | (~new_n365_ & ~new_n270_) | (~new_n247_ & ~new_n358_ & DATAI_22_) | ((new_n370_ | new_n247_) & new_n270_ & (~new_n247_ | new_n358_ | ~DATAI_22_))) & ((~new_n374_ & new_n247_ & new_n270_) | (~new_n247_ & ~new_n358_ & DATAI_23_) | (~new_n370_ & ~new_n270_) | ((new_n374_ | new_n247_) & new_n270_ & (~new_n247_ | new_n358_ | ~DATAI_23_)));
  assign new_n374_ = new_n376_ & (~new_n366_ | ~new_n375_);
  assign new_n375_ = REG3_REG_23__SCAN_IN ^ (REG3_REG_22__SCAN_IN & REG3_REG_21__SCAN_IN & REG3_REG_20__SCAN_IN & REG3_REG_19__SCAN_IN & new_n355_ & REG3_REG_18__SCAN_IN);
  assign new_n376_ = (~REG2_REG_23__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG0_REG_23__SCAN_IN | ~new_n254_ | new_n257_) & (~REG1_REG_23__SCAN_IN | new_n254_ | new_n257_);
  assign new_n377_ = (((new_n374_ | ~new_n247_ | ~new_n270_) & (new_n370_ | new_n270_) & (new_n247_ | ~new_n381_)) | (~new_n374_ & ~new_n247_) | ~new_n270_ | (new_n247_ & new_n381_)) & ((~new_n378_ & ~new_n247_) | ~new_n270_ | (new_n247_ & new_n382_) | ((new_n378_ | ~new_n247_ | ~new_n270_) & (new_n374_ | new_n270_) & (new_n247_ | ~new_n382_)));
  assign new_n378_ = new_n380_ & ((~new_n379_ & ~REG3_REG_24__SCAN_IN) | ~new_n366_ | (new_n379_ & REG3_REG_24__SCAN_IN));
  assign new_n379_ = REG3_REG_23__SCAN_IN & REG3_REG_22__SCAN_IN & REG3_REG_21__SCAN_IN & REG3_REG_20__SCAN_IN & REG3_REG_19__SCAN_IN & new_n355_ & REG3_REG_18__SCAN_IN;
  assign new_n380_ = (~REG1_REG_24__SCAN_IN | new_n254_ | new_n257_) & (~REG0_REG_24__SCAN_IN | ~new_n254_ | new_n257_) & (~REG2_REG_24__SCAN_IN | ~new_n254_ | ~new_n257_);
  assign new_n381_ = DATAI_23_ & (~new_n262_ | new_n265_ | (new_n263_ & ~new_n264_));
  assign new_n382_ = DATAI_24_ & (~new_n262_ | new_n265_ | (new_n263_ & ~new_n264_));
  assign new_n383_ = (((new_n348_ | ~new_n247_ | ~new_n270_) & (new_n247_ | new_n350_) & (new_n344_ | new_n270_)) | ~new_n270_ | (new_n247_ & ~new_n350_) | (~new_n247_ & ~new_n348_)) & (~new_n270_ | (new_n247_ & ~new_n384_) | (~new_n247_ & ~new_n359_) | ((new_n359_ | ~new_n247_ | ~new_n270_) & (new_n348_ | new_n270_) & (new_n247_ | new_n384_)));
  assign new_n384_ = (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) ? new_n385_ : ~DATAI_18_;
  assign new_n385_ = ((IR_REG_18__SCAN_IN & (~new_n363_ | ~new_n249_ | ~new_n250_)) | ~IR_REG_31__SCAN_IN | (~IR_REG_18__SCAN_IN & new_n363_ & new_n249_ & new_n250_)) & (~IR_REG_18__SCAN_IN | IR_REG_31__SCAN_IN);
  assign new_n386_ = ((~new_n359_ & new_n247_ & new_n270_) | (~new_n247_ & ~new_n384_) | (~new_n348_ & ~new_n270_) | (new_n270_ & (~new_n247_ | new_n384_) & (new_n247_ | new_n359_))) & ((new_n270_ & (~new_n247_ | new_n361_) & (new_n247_ | new_n360_)) | (~new_n360_ & new_n247_ & new_n270_) | (~new_n359_ & ~new_n270_) | (~new_n247_ & ~new_n361_));
  assign new_n387_ = ~new_n388_ & (((new_n392_ | new_n270_) & (new_n247_ | ~new_n397_) & (new_n395_ | ~new_n247_ | ~new_n270_)) | (~new_n395_ & ~new_n247_) | ~new_n270_ | (new_n247_ & new_n397_));
  assign new_n388_ = ((~new_n390_ & new_n270_ & new_n248_ & new_n252_) | (new_n389_ & (~new_n248_ | ~new_n252_))) & (new_n248_ | new_n390_ | new_n391_) & (new_n390_ | new_n252_) & (~new_n389_ | ~new_n270_ | ~new_n248_ | ~new_n252_);
  assign new_n389_ = ~new_n358_ & DATAI_30_;
  assign new_n390_ = (~REG0_REG_30__SCAN_IN | ~new_n254_ | new_n257_) & (~REG2_REG_30__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG1_REG_30__SCAN_IN | new_n254_ | new_n257_);
  assign new_n391_ = (~REG2_REG_31__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG0_REG_31__SCAN_IN | ~new_n254_ | new_n257_) & (~REG1_REG_31__SCAN_IN | new_n254_ | new_n257_);
  assign new_n392_ = new_n394_ & (~new_n366_ | (~REG3_REG_28__SCAN_IN & (~REG3_REG_27__SCAN_IN | ~REG3_REG_26__SCAN_IN | ~new_n393_ | ~REG3_REG_25__SCAN_IN)) | (REG3_REG_28__SCAN_IN & REG3_REG_27__SCAN_IN & REG3_REG_26__SCAN_IN & new_n393_ & REG3_REG_25__SCAN_IN));
  assign new_n393_ = REG3_REG_24__SCAN_IN & REG3_REG_23__SCAN_IN & REG3_REG_22__SCAN_IN & REG3_REG_21__SCAN_IN & REG3_REG_20__SCAN_IN & REG3_REG_19__SCAN_IN & new_n355_ & REG3_REG_18__SCAN_IN;
  assign new_n394_ = (~REG0_REG_28__SCAN_IN | ~new_n254_ | new_n257_) & (~REG2_REG_28__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG1_REG_28__SCAN_IN | new_n254_ | new_n257_);
  assign new_n395_ = new_n396_ & (~new_n366_ | ~REG3_REG_28__SCAN_IN | ~REG3_REG_27__SCAN_IN | ~REG3_REG_26__SCAN_IN | ~new_n393_ | ~REG3_REG_25__SCAN_IN);
  assign new_n396_ = (~REG0_REG_29__SCAN_IN | ~new_n254_ | new_n257_) & (~REG2_REG_29__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG1_REG_29__SCAN_IN | new_n254_ | new_n257_);
  assign new_n397_ = DATAI_29_ & (~new_n262_ | new_n265_ | (new_n263_ & ~new_n264_));
  assign new_n398_ = ((~new_n378_ & new_n247_ & new_n270_) | (~new_n374_ & ~new_n270_) | (~new_n247_ & new_n382_) | ((new_n378_ | new_n247_) & new_n270_ & (~new_n247_ | ~new_n382_))) & (((new_n399_ | new_n247_) & new_n270_ & (~new_n247_ | ~new_n401_)) | (~new_n399_ & new_n247_ & new_n270_) | (~new_n378_ & ~new_n270_) | (~new_n247_ & new_n401_));
  assign new_n399_ = new_n400_ & ((~new_n393_ & ~REG3_REG_25__SCAN_IN) | ~new_n366_ | (new_n393_ & REG3_REG_25__SCAN_IN));
  assign new_n400_ = (~REG1_REG_25__SCAN_IN | new_n254_ | new_n257_) & (~REG0_REG_25__SCAN_IN | ~new_n254_ | new_n257_) & (~REG2_REG_25__SCAN_IN | ~new_n254_ | ~new_n257_);
  assign new_n401_ = DATAI_25_ & (~new_n262_ | new_n265_ | (new_n263_ & ~new_n264_));
  assign new_n402_ = (((new_n399_ | ~new_n247_ | ~new_n270_) & (new_n378_ | new_n270_) & (new_n247_ | ~new_n401_)) | (~new_n399_ & ~new_n247_) | ~new_n270_ | (new_n247_ & new_n401_)) & (((new_n403_ | ~new_n247_ | ~new_n270_) & (~new_n405_ | new_n247_) & (new_n399_ | new_n270_)) | (~new_n403_ & ~new_n247_) | ~new_n270_ | (new_n405_ & new_n247_));
  assign new_n403_ = new_n404_ & (~new_n366_ | (REG3_REG_26__SCAN_IN & new_n393_ & REG3_REG_25__SCAN_IN) | (~REG3_REG_26__SCAN_IN & (~new_n393_ | ~REG3_REG_25__SCAN_IN)));
  assign new_n404_ = (~REG2_REG_26__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG0_REG_26__SCAN_IN | ~new_n254_ | new_n257_) & (~REG1_REG_26__SCAN_IN | new_n254_ | new_n257_);
  assign new_n405_ = ~new_n358_ & DATAI_26_;
  assign new_n406_ = ((~new_n403_ & new_n247_ & new_n270_) | (new_n405_ & ~new_n247_) | (~new_n399_ & ~new_n270_) | ((new_n403_ | new_n247_) & new_n270_ & (~new_n405_ | ~new_n247_))) & ((~new_n407_ & new_n247_ & new_n270_) | (~new_n403_ & ~new_n270_) | (new_n409_ & ~new_n247_) | (new_n270_ & (~new_n409_ | ~new_n247_) & (new_n407_ | new_n247_)));
  assign new_n407_ = new_n408_ & ((~REG3_REG_27__SCAN_IN & (~REG3_REG_26__SCAN_IN | ~new_n393_ | ~REG3_REG_25__SCAN_IN)) | ~new_n366_ | (REG3_REG_27__SCAN_IN & REG3_REG_26__SCAN_IN & new_n393_ & REG3_REG_25__SCAN_IN));
  assign new_n408_ = (~REG0_REG_27__SCAN_IN | ~new_n254_ | new_n257_) & (~REG2_REG_27__SCAN_IN | ~new_n254_ | ~new_n257_) & (~REG1_REG_27__SCAN_IN | new_n254_ | new_n257_);
  assign new_n409_ = ~new_n358_ & DATAI_27_;
  assign new_n410_ = (((new_n407_ | ~new_n247_ | ~new_n270_) & (new_n403_ | new_n270_) & (~new_n409_ | new_n247_)) | (~new_n407_ & ~new_n247_) | ~new_n270_ | (new_n409_ & new_n247_)) & (((new_n392_ | ~new_n247_ | ~new_n270_) & (new_n407_ | new_n270_) & (new_n247_ | ~new_n411_)) | (~new_n392_ & ~new_n247_) | ~new_n270_ | (new_n247_ & new_n411_));
  assign new_n411_ = DATAI_28_ & (~new_n262_ | new_n265_ | (new_n263_ & ~new_n264_));
  assign new_n412_ = ((~new_n392_ & new_n247_ & new_n270_) | (~new_n407_ & ~new_n270_) | (~new_n247_ & new_n411_) | ((new_n392_ | new_n247_) & new_n270_ & (~new_n247_ | ~new_n411_))) & (((new_n395_ | new_n247_) & new_n270_ & (~new_n247_ | ~new_n397_)) | (~new_n392_ & ~new_n270_) | (~new_n247_ & new_n397_) | (~new_n395_ & new_n247_ & new_n270_));
  assign new_n413_ = ((~new_n390_ & new_n270_ & new_n248_ & new_n252_) | ((~new_n248_ | ~new_n252_) & ~new_n358_ & DATAI_30_) | ((new_n248_ | new_n390_ | new_n391_) & (new_n390_ | new_n252_) & (~new_n270_ | ~new_n248_ | ~new_n252_ | new_n358_ | ~DATAI_30_))) & ((~new_n270_ & new_n248_ & new_n252_) | (~new_n391_ ^ (new_n358_ | ~DATAI_31_)));
  assign new_n414_ = (~new_n450_ | (~new_n415_ & new_n435_)) & new_n460_ & new_n453_ & (new_n439_ | ~new_n448_);
  assign new_n415_ = ~new_n433_ & ((new_n392_ & new_n411_) | (new_n416_ & (~new_n431_ | (new_n434_ & new_n418_ & new_n422_))));
  assign new_n416_ = ~new_n417_ & (new_n407_ | new_n409_);
  assign new_n417_ = ~new_n411_ & (~new_n394_ | (new_n366_ & (REG3_REG_28__SCAN_IN | (REG3_REG_27__SCAN_IN & REG3_REG_26__SCAN_IN & new_n393_ & REG3_REG_25__SCAN_IN)) & (~REG3_REG_28__SCAN_IN | ~REG3_REG_27__SCAN_IN | ~REG3_REG_26__SCAN_IN | ~new_n393_ | ~REG3_REG_25__SCAN_IN)));
  assign new_n418_ = new_n419_ & ~new_n420_ & ~new_n421_;
  assign new_n419_ = (new_n401_ | (new_n400_ & ((~REG3_REG_25__SCAN_IN & (~new_n379_ | ~REG3_REG_24__SCAN_IN)) | ~new_n366_ | (REG3_REG_25__SCAN_IN & new_n379_ & REG3_REG_24__SCAN_IN)))) & (new_n382_ | (new_n380_ & ((~new_n379_ & ~REG3_REG_24__SCAN_IN) | ~new_n366_ | (new_n379_ & REG3_REG_24__SCAN_IN))));
  assign new_n420_ = (~new_n382_ | ~new_n380_ | ((new_n379_ | REG3_REG_24__SCAN_IN) & new_n366_ & (~new_n379_ | ~REG3_REG_24__SCAN_IN))) & ~new_n381_ & (~new_n376_ | (new_n366_ & new_n375_));
  assign new_n421_ = (~new_n404_ | (new_n366_ & (~REG3_REG_26__SCAN_IN | ~new_n393_ | ~REG3_REG_25__SCAN_IN) & (REG3_REG_26__SCAN_IN | (new_n393_ & REG3_REG_25__SCAN_IN)))) & (new_n358_ | ~DATAI_26_);
  assign new_n422_ = (~new_n424_ | new_n423_ | new_n425_) & new_n428_ & ~new_n426_ & ~new_n427_ & new_n429_ & new_n430_;
  assign new_n423_ = new_n382_ & new_n380_ & ((~new_n379_ & ~REG3_REG_24__SCAN_IN) | ~new_n366_ | (new_n379_ & REG3_REG_24__SCAN_IN));
  assign new_n424_ = (new_n358_ | ~DATAI_22_) & (~new_n372_ | ((new_n371_ | REG3_REG_22__SCAN_IN) & new_n366_ & (~new_n371_ | ~REG3_REG_22__SCAN_IN)));
  assign new_n425_ = new_n381_ & new_n376_ & (~new_n366_ | ~new_n375_);
  assign new_n426_ = ~new_n368_ & (~new_n367_ | ((REG3_REG_21__SCAN_IN | (REG3_REG_20__SCAN_IN & REG3_REG_19__SCAN_IN & new_n355_ & REG3_REG_18__SCAN_IN)) & new_n366_ & (~REG3_REG_21__SCAN_IN | ~REG3_REG_20__SCAN_IN | ~REG3_REG_19__SCAN_IN | ~new_n355_ | ~REG3_REG_18__SCAN_IN)));
  assign new_n427_ = (new_n358_ | ~DATAI_20_) & (new_n354_ | ~new_n356_);
  assign new_n428_ = (new_n344_ | ~new_n345_) & (new_n359_ | ~new_n384_) & (new_n360_ | ~new_n361_) & (new_n348_ | ~new_n350_ | (new_n359_ & ~new_n384_));
  assign new_n429_ = (~new_n318_ | new_n322_) & (new_n320_ | new_n325_);
  assign new_n430_ = (new_n335_ | ~new_n336_) & (new_n339_ | ~new_n341_);
  assign new_n431_ = ~new_n432_ & (~new_n407_ | ~new_n409_) & (new_n421_ | ~new_n399_ | ~new_n401_);
  assign new_n432_ = new_n404_ & (~new_n366_ | (REG3_REG_26__SCAN_IN & new_n393_ & REG3_REG_25__SCAN_IN) | (~REG3_REG_26__SCAN_IN & (~new_n393_ | ~REG3_REG_25__SCAN_IN))) & ~new_n358_ & DATAI_26_;
  assign new_n433_ = ~new_n397_ & (~new_n396_ | (new_n366_ & REG3_REG_28__SCAN_IN & REG3_REG_27__SCAN_IN & REG3_REG_26__SCAN_IN & new_n393_ & REG3_REG_25__SCAN_IN));
  assign new_n434_ = new_n327_ & ~new_n329_;
  assign new_n435_ = (~new_n436_ | ~new_n418_ | ~new_n422_) & (~new_n389_ | ~new_n390_) & (~new_n395_ | ~new_n397_);
  assign new_n436_ = ~new_n417_ & (new_n407_ | new_n409_) & ~new_n433_ & ~new_n437_ & new_n438_;
  assign new_n437_ = ((~new_n306_ & ~new_n310_) | (~new_n301_ & new_n307_) | ((new_n287_ | ~new_n291_) & (~new_n306_ | ~new_n310_))) & (~new_n299_ | new_n303_) & (~new_n301_ | new_n307_);
  assign new_n438_ = (new_n299_ | ~new_n303_) & ((new_n320_ & new_n325_) | new_n327_ | ~new_n329_);
  assign new_n439_ = (new_n440_ | ~new_n441_ | new_n447_ | (~new_n283_ & new_n284_ & (~new_n289_ | ~new_n293_))) & (~new_n441_ | ~new_n442_) & (new_n440_ | ~new_n441_ | ~new_n283_ | new_n284_);
  assign new_n440_ = new_n424_ & ~new_n423_ & ~new_n425_;
  assign new_n441_ = new_n429_ & new_n430_ & new_n428_ & ~new_n426_ & ~new_n427_;
  assign new_n442_ = ~new_n424_ & new_n444_ & new_n443_ & ~new_n445_ & (new_n283_ | ~new_n284_ | (new_n289_ & new_n293_));
  assign new_n443_ = (new_n253_ | ~new_n261_) & (new_n260_ | ~new_n268_);
  assign new_n444_ = (new_n272_ | ~new_n277_) & (new_n267_ | new_n273_) & (~new_n275_ | new_n276_);
  assign new_n445_ = (new_n275_ | ~new_n276_) & new_n446_ & (new_n252_ | ~new_n362_);
  assign new_n446_ = IR_REG_21__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_20__SCAN_IN & new_n251_ & new_n249_ & new_n250_));
  assign new_n447_ = (~new_n253_ | new_n261_) & ((~new_n260_ & new_n268_) | (~new_n253_ & new_n261_) | ((~new_n272_ | new_n277_ | (~new_n267_ & ~new_n273_)) & (~new_n267_ | ~new_n273_) & (~new_n260_ | new_n268_)));
  assign new_n448_ = new_n449_ & (new_n289_ | new_n293_) & new_n451_ & new_n452_;
  assign new_n449_ = ~new_n417_ & (new_n407_ | new_n409_) & new_n450_ & ~new_n433_ & new_n419_ & ~new_n420_ & ~new_n421_;
  assign new_n450_ = (~new_n391_ | new_n358_ | ~DATAI_31_) & (new_n390_ | (~new_n358_ & DATAI_30_));
  assign new_n451_ = (new_n301_ | ~new_n307_) & (new_n306_ | new_n310_);
  assign new_n452_ = ((new_n320_ & new_n325_) | new_n327_ | ~new_n329_) & (new_n299_ | ~new_n303_) & (~new_n287_ | new_n291_);
  assign new_n453_ = ~new_n458_ & (new_n440_ | ~new_n449_ | (new_n454_ & (~new_n441_ | ~new_n457_) & (new_n426_ | ~new_n459_)));
  assign new_n454_ = ~new_n423_ & ~new_n425_ & ~new_n455_ & ~new_n456_;
  assign new_n455_ = ~new_n358_ & DATAI_22_ & new_n372_ & ((~new_n371_ & ~REG3_REG_22__SCAN_IN) | ~new_n366_ | (new_n371_ & REG3_REG_22__SCAN_IN));
  assign new_n456_ = new_n368_ & new_n367_ & ((~REG3_REG_21__SCAN_IN & (~REG3_REG_20__SCAN_IN | ~REG3_REG_19__SCAN_IN | ~new_n355_ | ~REG3_REG_18__SCAN_IN)) | ~new_n366_ | (REG3_REG_21__SCAN_IN & REG3_REG_20__SCAN_IN & REG3_REG_19__SCAN_IN & new_n355_ & REG3_REG_18__SCAN_IN));
  assign new_n457_ = new_n451_ & new_n452_ & new_n289_ & new_n293_;
  assign new_n458_ = ~new_n391_ & (new_n358_ | ~DATAI_31_);
  assign new_n459_ = ~new_n358_ & DATAI_20_ & ~new_n354_ & new_n356_;
  assign new_n460_ = (~new_n462_ | ~new_n461_ | new_n440_ | ~new_n449_) & (new_n465_ | ~new_n461_ | new_n440_ | ~new_n449_) & (new_n466_ | new_n440_ | ~new_n449_ | ~new_n461_ | ~new_n428_) & (~new_n464_ | new_n440_ | ~new_n449_ | ~new_n461_ | ~new_n428_);
  assign new_n461_ = ~new_n426_ & ~new_n427_;
  assign new_n462_ = new_n463_ & (new_n360_ | ~new_n361_);
  assign new_n463_ = new_n359_ & ~new_n384_;
  assign new_n464_ = new_n430_ & new_n320_ & new_n325_ & (~new_n318_ | new_n322_);
  assign new_n465_ = (~new_n360_ | new_n361_) & ((~new_n359_ & new_n384_) | (~new_n360_ & new_n361_) | ((~new_n348_ | new_n350_) & (~new_n344_ | new_n345_ | (~new_n348_ & new_n350_ & (~new_n359_ | new_n384_)))));
  assign new_n466_ = (new_n318_ | ~new_n322_ | (~new_n335_ & new_n336_) | (~new_n339_ & new_n341_)) & (~new_n339_ | new_n341_) & (~new_n335_ | new_n336_ | (~new_n339_ & new_n341_));
  assign new_n467_ = new_n488_ & new_n492_ & new_n493_ & new_n489_ & (new_n490_ | new_n491_) & new_n468_ & new_n470_;
  assign new_n468_ = ~new_n469_ & ~new_n423_;
  assign new_n469_ = ~new_n378_ & ~new_n382_;
  assign new_n470_ = new_n486_ & new_n484_ & new_n485_ & new_n479_ & new_n473_ & new_n476_ & new_n471_ & ~new_n427_;
  assign new_n471_ = ~new_n472_ & (new_n360_ | ~new_n361_);
  assign new_n472_ = ~new_n359_ & new_n384_;
  assign new_n473_ = new_n475_ & new_n474_ & (new_n272_ | ~new_n277_) & (~new_n272_ | new_n277_) & (new_n287_ ^ ~new_n291_);
  assign new_n474_ = (new_n299_ | ~new_n303_) & (new_n327_ | ~new_n329_) & (new_n260_ | ~new_n268_) & (~new_n260_ | new_n268_);
  assign new_n475_ = (~new_n339_ | new_n341_) & (new_n339_ | ~new_n341_) & (new_n289_ ^ new_n293_) & (~new_n299_ | new_n303_) & (~new_n301_ | new_n307_);
  assign new_n476_ = (new_n344_ ^ ~new_n345_) & new_n478_ & new_n477_ & (new_n267_ ^ new_n273_);
  assign new_n477_ = ~new_n318_ ^ new_n322_;
  assign new_n478_ = (new_n253_ | ~new_n261_) & (~new_n253_ | new_n261_) & (~new_n320_ | ~new_n325_) & (~new_n327_ | new_n329_);
  assign new_n479_ = (new_n348_ | ~new_n350_) & (~new_n348_ | new_n350_) & ~new_n463_ & new_n482_ & new_n483_ & new_n480_ & new_n481_;
  assign new_n480_ = (~new_n275_ | new_n276_) & (new_n275_ | ~new_n276_) & (new_n320_ | new_n325_) & (new_n390_ | (~new_n358_ & DATAI_30_));
  assign new_n481_ = (new_n391_ | (~new_n358_ & DATAI_31_)) & (~new_n391_ | new_n358_ | ~DATAI_31_) & (new_n306_ | new_n310_) & (new_n301_ | ~new_n307_);
  assign new_n482_ = ~new_n335_ ^ new_n336_;
  assign new_n483_ = (~new_n283_ | new_n284_) & (new_n283_ | ~new_n284_) & (~new_n306_ | ~new_n310_) & (~new_n390_ | new_n358_ | ~DATAI_30_);
  assign new_n484_ = ~new_n459_ & (~new_n360_ | new_n361_);
  assign new_n485_ = ~new_n426_ & ~new_n456_;
  assign new_n486_ = ~new_n487_ & ~new_n425_ & ~new_n424_ & ~new_n455_;
  assign new_n487_ = ~new_n381_ & (~new_n376_ | (new_n366_ & new_n375_));
  assign new_n488_ = ~new_n392_ ^ (new_n358_ | ~DATAI_28_);
  assign new_n489_ = ~new_n421_ & ~new_n432_;
  assign new_n490_ = new_n399_ & ~new_n401_;
  assign new_n491_ = ~new_n399_ & new_n401_;
  assign new_n492_ = ~new_n395_ ^ (new_n358_ | ~DATAI_29_);
  assign new_n493_ = ~new_n407_ ^ ~new_n409_;
  assign new_n494_ = ((new_n247_ & new_n270_) | (~new_n391_ & (new_n358_ | ~DATAI_31_))) & (~new_n247_ | (new_n391_ & ~new_n358_ & DATAI_31_));
  assign new_n495_ = new_n496_ & (~new_n525_ | new_n242_ | new_n494_);
  assign new_n496_ = ~new_n497_ & ~new_n523_ & (~new_n414_ | ((~new_n248_ | new_n446_ | ~new_n362_) & (~new_n362_ | ~new_n248_ | ~new_n252_))) & (new_n467_ | ~new_n362_ | new_n248_ | ~new_n446_);
  assign new_n497_ = new_n522_ & new_n521_ & (~new_n517_ | (new_n520_ & (~new_n515_ | (new_n419_ & (new_n498_ | ~new_n519_)))));
  assign new_n498_ = new_n500_ & (~new_n499_ | (~new_n427_ & (~new_n514_ | (new_n512_ & (~new_n510_ | (~new_n501_ & new_n509_))))));
  assign new_n499_ = ~new_n455_ & ~new_n456_;
  assign new_n500_ = (~new_n426_ | new_n455_) & ~new_n487_ & ~new_n424_;
  assign new_n501_ = new_n503_ & (~new_n451_ | (new_n502_ & (new_n505_ | ~new_n508_ | (new_n507_ & ~new_n504_ & ~new_n506_))));
  assign new_n502_ = (new_n287_ | ~new_n291_) & (~new_n306_ | ~new_n310_);
  assign new_n503_ = (~new_n299_ | new_n303_) & (~new_n301_ | new_n307_);
  assign new_n504_ = new_n253_ & ~new_n261_;
  assign new_n505_ = new_n287_ & ~new_n291_;
  assign new_n506_ = (new_n260_ | ~new_n268_) & ((new_n260_ & ~new_n268_) | (new_n267_ & new_n273_) | ((new_n267_ | new_n273_) & ((new_n272_ & ~new_n277_) | (~new_n275_ & new_n276_ & (new_n272_ | ~new_n277_)))));
  assign new_n507_ = (~new_n283_ | new_n284_) & (~new_n289_ | ~new_n293_);
  assign new_n508_ = (new_n289_ | new_n293_) & (((new_n253_ | ~new_n261_) & (new_n283_ | ~new_n284_)) | (new_n283_ & ~new_n284_) | (new_n289_ & new_n293_));
  assign new_n509_ = new_n429_ & (new_n299_ | ~new_n303_) & (new_n327_ | ~new_n329_);
  assign new_n510_ = new_n511_ & (~new_n434_ | (~new_n320_ & ~new_n325_) | (new_n318_ & ~new_n322_)) & (new_n318_ | ~new_n322_) & (~new_n320_ | ~new_n325_ | (new_n318_ & ~new_n322_));
  assign new_n511_ = (~new_n335_ | new_n336_) & (~new_n339_ | new_n341_) & (~new_n344_ | new_n345_);
  assign new_n512_ = new_n513_ & (new_n344_ | ~new_n345_) & ~new_n472_ & (new_n360_ | ~new_n361_);
  assign new_n513_ = (new_n348_ | ~new_n350_) & (((new_n335_ | ~new_n336_) & (new_n339_ | ~new_n341_)) | (new_n339_ & ~new_n341_) | (new_n344_ & ~new_n345_));
  assign new_n514_ = ~new_n459_ & (~new_n360_ | new_n361_) & ((~new_n360_ & new_n361_) | (~new_n359_ & new_n384_) | ((~new_n359_ | new_n384_) & (~new_n348_ | new_n350_)));
  assign new_n515_ = ~new_n516_ & ~new_n432_;
  assign new_n516_ = new_n399_ & new_n401_;
  assign new_n517_ = new_n518_ & (~new_n395_ | ~new_n397_) & (~new_n392_ | ~new_n411_) & (~new_n407_ | ~new_n409_);
  assign new_n518_ = ~new_n458_ & (~new_n389_ | (~new_n390_ & ~new_n391_));
  assign new_n519_ = ~new_n423_ & ~new_n425_;
  assign new_n520_ = ~new_n421_ & (new_n407_ | new_n409_);
  assign new_n521_ = (~new_n417_ | (new_n395_ & ~new_n358_ & DATAI_29_) | (~new_n391_ & (new_n358_ | ~DATAI_31_)) | ((new_n390_ | new_n391_) & ~new_n358_ & DATAI_30_)) & ((~new_n391_ & (new_n358_ | ~DATAI_31_)) | ((new_n390_ | new_n391_) & ~new_n358_ & DATAI_30_) | new_n395_ | (~new_n358_ & DATAI_29_)) & (new_n358_ | ~DATAI_31_ | (~new_n391_ & (new_n390_ | (~new_n358_ & DATAI_30_))));
  assign new_n522_ = ~new_n248_ & ~new_n446_ & ~new_n252_ & ~new_n362_;
  assign new_n523_ = new_n524_ & (~new_n521_ | (new_n517_ & (~new_n520_ | (new_n515_ & (~new_n419_ | (~new_n498_ & new_n519_))))));
  assign new_n524_ = new_n362_ & ~new_n248_ & ~new_n446_;
  assign new_n525_ = new_n362_ & new_n526_;
  assign new_n526_ = (~IR_REG_20__SCAN_IN | IR_REG_31__SCAN_IN) & ((IR_REG_20__SCAN_IN & (~new_n251_ | ~new_n249_ | ~new_n250_)) | ~IR_REG_31__SCAN_IN | (~IR_REG_20__SCAN_IN & new_n251_ & new_n249_ & new_n250_)) & (IR_REG_22__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (new_n251_ & new_n249_ & new_n250_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN))) & (~IR_REG_21__SCAN_IN | (IR_REG_31__SCAN_IN & (IR_REG_20__SCAN_IN | ~new_n251_ | ~new_n249_ | ~new_n250_))) & (IR_REG_21__SCAN_IN | ~IR_REG_31__SCAN_IN | (~IR_REG_20__SCAN_IN & new_n251_ & new_n249_ & new_n250_));
  assign new_n527_ = ~new_n583_ & new_n596_ & ((new_n582_ & (new_n528_ | new_n581_)) | ~new_n601_ | (~new_n528_ & ~new_n581_ & ~new_n582_));
  assign new_n528_ = new_n580_ & (~new_n575_ | (~new_n579_ & (new_n577_ | (new_n578_ ^ new_n536_)) & ((~new_n529_ & new_n573_) | (new_n577_ & (~new_n578_ | ~new_n536_) & (new_n578_ | new_n536_)))));
  assign new_n529_ = new_n568_ & new_n572_ & (~new_n565_ | (new_n563_ & (new_n569_ | (~new_n571_ & (new_n530_ | new_n570_)))));
  assign new_n530_ = ~new_n559_ & (~new_n555_ | (new_n551_ & ~new_n560_ & (new_n561_ | (~new_n562_ & (new_n531_ | ~new_n547_)))));
  assign new_n531_ = new_n532_ & new_n546_ & (new_n538_ | new_n545_ | (new_n544_ & ~new_n539_ & (new_n540_ | new_n541_)));
  assign new_n532_ = ((~new_n536_ & ((new_n293_ & new_n535_) | (~new_n289_ & new_n533_))) | (new_n536_ & (~new_n293_ | ~new_n535_) & (new_n289_ | ~new_n533_)) | (new_n293_ & new_n533_) | (~new_n289_ & new_n537_)) & ((~new_n536_ & ((~new_n287_ & new_n535_) | (~new_n291_ & new_n533_))) | (new_n536_ & (new_n287_ | ~new_n535_) & (new_n291_ | ~new_n533_)) | (~new_n287_ & new_n533_) | (~new_n291_ & new_n537_));
  assign new_n533_ = ~new_n534_ & new_n248_ & ~new_n446_;
  assign new_n534_ = ((IR_REG_26__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & (IR_REG_26__SCAN_IN | IR_REG_25__SCAN_IN | IR_REG_24__SCAN_IN | ~new_n249_ | ~new_n250_ | ~new_n251_ | ~new_n255_) & (~IR_REG_26__SCAN_IN | (~IR_REG_25__SCAN_IN & ~IR_REG_24__SCAN_IN & new_n249_ & new_n250_ & new_n251_ & new_n255_)))) & ((IR_REG_24__SCAN_IN & ~IR_REG_31__SCAN_IN) | ((~IR_REG_24__SCAN_IN | (new_n249_ & new_n250_ & new_n251_ & new_n255_)) & IR_REG_31__SCAN_IN & (IR_REG_24__SCAN_IN | ~new_n249_ | ~new_n250_ | ~new_n251_ | ~new_n255_))) & (~IR_REG_25__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_24__SCAN_IN & new_n249_ & new_n250_ & new_n251_ & new_n255_)));
  assign new_n535_ = ~new_n534_ & ((~new_n252_ & new_n446_) | ~new_n248_ | (new_n362_ ? new_n446_ : new_n252_));
  assign new_n536_ = ~new_n534_ & (~new_n248_ | new_n446_) & (new_n362_ | ~new_n252_ | ~new_n446_);
  assign new_n537_ = ~new_n534_ & (~new_n248_ | (new_n362_ ? new_n446_ : new_n252_));
  assign new_n538_ = ((~new_n253_ & new_n537_) | (~new_n261_ & new_n533_)) & (new_n536_ ^ ((~new_n253_ & new_n533_) | (~new_n261_ & new_n535_)));
  assign new_n539_ = (new_n272_ | ~new_n537_) & (new_n277_ | ~new_n533_) & (new_n536_ | ((new_n272_ | ~new_n533_) & (new_n277_ | ~new_n535_))) & (~new_n536_ | (~new_n272_ & new_n533_) | (~new_n277_ & new_n535_));
  assign new_n540_ = ((~new_n272_ & new_n537_) | (~new_n277_ & new_n533_)) & (new_n536_ ^ ((~new_n272_ & new_n533_) | (~new_n277_ & new_n535_)));
  assign new_n541_ = ((new_n276_ | ~new_n533_) & ~new_n542_ & (new_n275_ | ~new_n535_)) ? new_n536_ : ((~new_n276_ & new_n537_) | new_n543_ | (~new_n275_ & new_n533_));
  assign new_n542_ = new_n534_ & REG1_REG_0__SCAN_IN;
  assign new_n543_ = new_n534_ & IR_REG_0__SCAN_IN;
  assign new_n544_ = ((~new_n536_ & ((new_n273_ & new_n535_) | (~new_n267_ & new_n533_))) | (new_n536_ & (~new_n273_ | ~new_n535_) & (new_n267_ | ~new_n533_)) | (new_n273_ & new_n533_) | (~new_n267_ & new_n537_)) & ((~new_n260_ & new_n537_) | (~new_n268_ & new_n533_) | (~new_n536_ & ((~new_n260_ & new_n533_) | (~new_n268_ & new_n535_))) | (new_n536_ & (new_n260_ | ~new_n533_) & (new_n268_ | ~new_n535_)));
  assign new_n545_ = ((~new_n260_ & new_n537_) | (~new_n268_ & new_n533_) | (~new_n536_ & ((~new_n260_ & new_n533_) | (~new_n268_ & new_n535_))) | (new_n536_ & (new_n260_ | ~new_n533_) & (new_n268_ | ~new_n535_))) & ((((~new_n260_ & new_n537_) | (~new_n268_ & new_n533_)) & (new_n536_ ^ ((~new_n260_ & new_n533_) | (~new_n268_ & new_n535_)))) | ((new_n536_ ^ ((new_n273_ & new_n535_) | (~new_n267_ & new_n533_))) & ((new_n273_ & new_n533_) | (~new_n267_ & new_n537_))));
  assign new_n546_ = ((~new_n284_ & new_n533_) | (~new_n283_ & new_n537_) | (~new_n536_ & ((~new_n284_ & new_n535_) | (~new_n283_ & new_n533_))) | (new_n536_ & (new_n284_ | ~new_n535_) & (new_n283_ | ~new_n533_))) & ((~new_n253_ & new_n537_) | (~new_n261_ & new_n533_) | (~new_n536_ & ((~new_n253_ & new_n533_) | (~new_n261_ & new_n535_))) | (new_n536_ & (new_n253_ | ~new_n533_) & (new_n261_ | ~new_n535_)));
  assign new_n547_ = ~new_n549_ & new_n550_ & (~new_n532_ | ~new_n548_);
  assign new_n548_ = ((~new_n283_ & new_n537_) | (~new_n284_ & new_n533_)) & (new_n536_ ^ ((~new_n283_ & new_n533_) | (~new_n284_ & new_n535_)));
  assign new_n549_ = ((~new_n536_ & ((~new_n287_ & new_n535_) | (~new_n291_ & new_n533_))) | (new_n536_ & (new_n287_ | ~new_n535_) & (new_n291_ | ~new_n533_)) | (~new_n287_ & new_n533_) | (~new_n291_ & new_n537_)) & (new_n536_ ^ ((new_n293_ & new_n535_) | (~new_n289_ & new_n533_))) & ((new_n293_ & new_n533_) | (~new_n289_ & new_n537_));
  assign new_n550_ = ((~new_n536_ ^ ((~new_n287_ & new_n535_) | (~new_n291_ & new_n533_))) | ((new_n287_ | ~new_n533_) & (new_n291_ | ~new_n537_))) & ((~new_n536_ ^ ((new_n310_ & new_n535_) | (~new_n306_ & new_n533_))) | ((~new_n310_ | ~new_n533_) & (new_n306_ | ~new_n537_)));
  assign new_n551_ = ~new_n554_ & new_n552_ & ~new_n553_;
  assign new_n552_ = ((~new_n536_ & ((new_n325_ & new_n535_) | (~new_n320_ & new_n533_))) | (new_n536_ & (~new_n325_ | ~new_n535_) & (new_n320_ | ~new_n533_)) | (new_n325_ & new_n533_) | (~new_n320_ & new_n537_)) & ((~new_n536_ & ((~new_n318_ & new_n535_) | (~new_n322_ & new_n533_))) | (new_n536_ & (new_n318_ | ~new_n535_) & (new_n322_ | ~new_n533_)) | (~new_n318_ & new_n533_) | (~new_n322_ & new_n537_));
  assign new_n553_ = (new_n327_ | ~new_n537_) & (new_n329_ | ~new_n533_) & (new_n536_ | ((new_n327_ | ~new_n533_) & (new_n329_ | ~new_n535_))) & (~new_n536_ | (~new_n327_ & new_n533_) | (~new_n329_ & new_n535_));
  assign new_n554_ = (new_n299_ | ~new_n537_) & (new_n303_ | ~new_n533_) & (new_n536_ | ((new_n299_ | ~new_n533_) & (new_n303_ | ~new_n535_))) & (~new_n536_ | (~new_n299_ & new_n533_) | (~new_n303_ & new_n535_));
  assign new_n555_ = (~new_n556_ | ~new_n552_ | new_n553_) & ~new_n557_ & (~new_n552_ | new_n558_);
  assign new_n556_ = ((~new_n299_ & new_n537_) | (~new_n303_ & new_n533_)) & (new_n536_ ^ ((~new_n299_ & new_n533_) | (~new_n303_ & new_n535_)));
  assign new_n557_ = (new_n536_ ^ ((~new_n318_ & new_n535_) | (~new_n322_ & new_n533_))) & ((~new_n318_ & new_n533_) | (~new_n322_ & new_n537_));
  assign new_n558_ = ((~new_n536_ ^ ((new_n325_ & new_n535_) | (~new_n320_ & new_n533_))) | ((~new_n325_ | ~new_n533_) & (new_n320_ | ~new_n537_))) & (((new_n329_ | ~new_n533_) & (new_n327_ | ~new_n537_)) | (~new_n536_ ^ ((~new_n329_ & new_n535_) | (~new_n327_ & new_n533_))));
  assign new_n559_ = (new_n335_ | ~new_n537_) & (new_n336_ | ~new_n533_) & (new_n536_ | ((new_n335_ | ~new_n533_) & (new_n336_ | ~new_n535_))) & (~new_n536_ | (~new_n335_ & new_n533_) | (~new_n336_ & new_n535_));
  assign new_n560_ = (new_n301_ | ~new_n537_) & (new_n307_ | ~new_n533_) & (new_n536_ | ((new_n301_ | ~new_n533_) & (new_n307_ | ~new_n535_))) & (~new_n536_ | (~new_n301_ & new_n533_) | (~new_n307_ & new_n535_));
  assign new_n561_ = ((~new_n301_ & new_n537_) | (~new_n307_ & new_n533_)) & (new_n536_ ^ ((~new_n301_ & new_n533_) | (~new_n307_ & new_n535_)));
  assign new_n562_ = (new_n536_ | ((new_n306_ | ~new_n533_) & (~new_n310_ | ~new_n535_))) & (~new_n536_ | (~new_n306_ & new_n533_) | (new_n310_ & new_n535_)) & (new_n306_ | ~new_n537_) & (~new_n310_ | ~new_n533_);
  assign new_n563_ = ~new_n564_ & ((~new_n350_ & new_n533_) | (~new_n348_ & new_n537_) | (~new_n536_ & ((~new_n348_ & new_n533_) | (~new_n350_ & new_n535_))) | (new_n536_ & (new_n348_ | ~new_n533_) & (new_n350_ | ~new_n535_)));
  assign new_n564_ = (new_n344_ | ~new_n537_) & (new_n345_ | ~new_n533_) & (new_n536_ | ((new_n344_ | ~new_n533_) & (new_n345_ | ~new_n535_))) & (~new_n536_ | (~new_n344_ & new_n533_) | (~new_n345_ & new_n535_));
  assign new_n565_ = (~new_n566_ | ((new_n350_ | ~new_n533_) & (new_n348_ | ~new_n537_) & (new_n536_ | ((new_n350_ | ~new_n535_) & (new_n348_ | ~new_n533_))) & (~new_n536_ | (~new_n350_ & new_n535_) | (~new_n348_ & new_n533_)))) & ~new_n567_ & (((new_n350_ | ~new_n533_) & (new_n348_ | ~new_n537_)) | (~new_n536_ ^ ((~new_n350_ & new_n535_) | (~new_n348_ & new_n533_))));
  assign new_n566_ = ((~new_n344_ & new_n537_) | (~new_n345_ & new_n533_)) & (new_n536_ ^ ((~new_n344_ & new_n533_) | (~new_n345_ & new_n535_)));
  assign new_n567_ = ((~new_n359_ & new_n537_) | (~new_n384_ & new_n533_)) & (new_n536_ ^ ((~new_n359_ & new_n533_) | (~new_n384_ & new_n535_)));
  assign new_n568_ = ((~new_n536_ & ((new_n368_ & new_n535_) | (~new_n365_ & new_n533_))) | (new_n536_ & (~new_n368_ | ~new_n535_) & (new_n365_ | ~new_n533_)) | (new_n368_ & new_n533_) | (~new_n365_ & new_n537_)) & ((~new_n536_ & ((new_n357_ & new_n535_) | (~new_n353_ & new_n533_))) | (new_n536_ & (~new_n357_ | ~new_n535_) & (new_n353_ | ~new_n533_)) | (new_n357_ & new_n533_) | (~new_n353_ & new_n537_));
  assign new_n569_ = ((~new_n339_ & new_n537_) | (~new_n341_ & new_n533_)) & (new_n536_ ^ ((~new_n339_ & new_n533_) | (~new_n341_ & new_n535_)));
  assign new_n570_ = ((~new_n335_ & new_n537_) | (~new_n336_ & new_n533_)) & (new_n536_ ^ ((~new_n335_ & new_n533_) | (~new_n336_ & new_n535_)));
  assign new_n571_ = (new_n339_ | ~new_n537_) & (new_n341_ | ~new_n533_) & (new_n536_ | ((new_n339_ | ~new_n533_) & (new_n341_ | ~new_n535_))) & (~new_n536_ | (~new_n339_ & new_n533_) | (~new_n341_ & new_n535_));
  assign new_n572_ = ((~new_n361_ & new_n533_) | (~new_n360_ & new_n537_) | (~new_n536_ & ((~new_n361_ & new_n535_) | (~new_n360_ & new_n533_))) | (new_n536_ & (new_n361_ | ~new_n535_) & (new_n360_ | ~new_n533_))) & ((~new_n359_ & new_n537_) | (~new_n384_ & new_n533_) | (~new_n536_ & ((~new_n359_ & new_n533_) | (~new_n384_ & new_n535_))) | (new_n536_ & (new_n359_ | ~new_n533_) & (new_n384_ | ~new_n535_)));
  assign new_n573_ = (~new_n568_ | new_n574_) & ((~new_n536_ ^ ((new_n368_ & new_n535_) | (~new_n365_ & new_n533_))) | ((~new_n368_ | ~new_n533_) & (new_n365_ | ~new_n537_)));
  assign new_n574_ = ((~new_n536_ ^ ((new_n357_ & new_n535_) | (~new_n353_ & new_n533_))) | ((~new_n357_ | ~new_n533_) & (new_n353_ | ~new_n537_))) & (((new_n361_ | ~new_n533_) & (new_n360_ | ~new_n537_)) | (~new_n536_ ^ ((~new_n361_ & new_n535_) | (~new_n360_ & new_n533_))));
  assign new_n575_ = ~new_n576_ & ((new_n382_ & new_n533_) | (~new_n378_ & new_n537_) | (~new_n536_ & ((new_n382_ & new_n535_) | (~new_n378_ & new_n533_))) | (new_n536_ & (~new_n382_ | ~new_n535_) & (new_n378_ | ~new_n533_)));
  assign new_n576_ = (new_n536_ | ((new_n374_ | ~new_n533_) & (~new_n381_ | ~new_n535_))) & (~new_n536_ | (~new_n374_ & new_n533_) | (new_n381_ & new_n535_)) & (new_n374_ | ~new_n537_) & (~new_n381_ | ~new_n533_);
  assign new_n577_ = (new_n370_ | ~new_n537_) & (~new_n533_ | new_n358_ | ~DATAI_22_);
  assign new_n578_ = (new_n370_ | ~new_n533_) & (~new_n535_ | new_n358_ | ~DATAI_22_);
  assign new_n579_ = (new_n536_ ^ ((~new_n374_ & new_n533_) | (new_n381_ & new_n535_))) & ((~new_n374_ & new_n537_) | (new_n381_ & new_n533_));
  assign new_n580_ = ((~new_n536_ ^ ((new_n401_ & new_n535_) | (~new_n399_ & new_n533_))) | ((~new_n401_ | ~new_n533_) & (new_n399_ | ~new_n537_))) & (((~new_n382_ | ~new_n533_) & (new_n378_ | ~new_n537_)) | (~new_n536_ ^ ((new_n382_ & new_n535_) | (~new_n378_ & new_n533_))));
  assign new_n581_ = (new_n536_ | ((new_n399_ | ~new_n533_) & (~new_n401_ | ~new_n535_))) & (~new_n536_ | (~new_n399_ & new_n533_) | (new_n401_ & new_n535_)) & (new_n399_ | ~new_n537_) & (~new_n401_ | ~new_n533_);
  assign new_n582_ = ((new_n403_ | ~new_n537_) & (~new_n405_ | ~new_n533_)) ^ (~new_n536_ ^ ((new_n403_ | ~new_n533_) & (~new_n405_ | ~new_n535_)));
  assign new_n583_ = new_n593_ & ((~new_n407_ & new_n584_ & new_n262_) | (~new_n399_ & new_n584_ & ~new_n262_) | (~new_n584_ & (~REG3_REG_26__SCAN_IN | ~new_n393_ | ~REG3_REG_25__SCAN_IN) & (REG3_REG_26__SCAN_IN | (new_n393_ & REG3_REG_25__SCAN_IN))));
  assign new_n584_ = (~new_n585_ | ~new_n587_) & (D_REG_1__SCAN_IN | (new_n587_ & new_n586_ & B_REG_SCAN_IN) | new_n585_ | (~new_n586_ & ~B_REG_SCAN_IN)) & (new_n588_ | (new_n587_ & new_n586_ & B_REG_SCAN_IN) | new_n585_ | (~new_n586_ & ~B_REG_SCAN_IN)) & (~new_n585_ | ~new_n586_) & (D_REG_0__SCAN_IN | (new_n587_ & new_n586_ & B_REG_SCAN_IN) | new_n585_ | (~new_n586_ & ~B_REG_SCAN_IN));
  assign new_n585_ = (~IR_REG_26__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_26__SCAN_IN & ~IR_REG_25__SCAN_IN & ~IR_REG_24__SCAN_IN & new_n249_ & new_n250_ & new_n251_ & new_n255_) | (IR_REG_26__SCAN_IN & (IR_REG_25__SCAN_IN | IR_REG_24__SCAN_IN | ~new_n249_ | ~new_n250_ | ~new_n251_ | ~new_n255_)));
  assign new_n586_ = (~IR_REG_24__SCAN_IN | IR_REG_31__SCAN_IN) & ((IR_REG_24__SCAN_IN & (~new_n249_ | ~new_n250_ | ~new_n251_ | ~new_n255_)) | ~IR_REG_31__SCAN_IN | (~IR_REG_24__SCAN_IN & new_n249_ & new_n250_ & new_n251_ & new_n255_));
  assign new_n587_ = IR_REG_25__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_24__SCAN_IN & new_n249_ & new_n250_ & new_n251_ & new_n255_));
  assign new_n588_ = new_n589_ & new_n590_ & new_n591_ & new_n592_;
  assign new_n589_ = ~D_REG_16__SCAN_IN & ~D_REG_17__SCAN_IN & ~D_REG_18__SCAN_IN & ~D_REG_19__SCAN_IN & ~D_REG_20__SCAN_IN & ~D_REG_21__SCAN_IN & ~D_REG_22__SCAN_IN & ~D_REG_23__SCAN_IN;
  assign new_n590_ = ~D_REG_24__SCAN_IN & ~D_REG_25__SCAN_IN & ~D_REG_26__SCAN_IN & ~D_REG_27__SCAN_IN & ~D_REG_28__SCAN_IN & ~D_REG_29__SCAN_IN & ~D_REG_30__SCAN_IN & ~D_REG_31__SCAN_IN;
  assign new_n591_ = ~D_REG_2__SCAN_IN & ~D_REG_3__SCAN_IN & ~D_REG_6__SCAN_IN & ~D_REG_7__SCAN_IN & ~D_REG_4__SCAN_IN & ~D_REG_5__SCAN_IN;
  assign new_n592_ = ~D_REG_8__SCAN_IN & ~D_REG_9__SCAN_IN & ~D_REG_10__SCAN_IN & ~D_REG_11__SCAN_IN & ~D_REG_12__SCAN_IN & ~D_REG_13__SCAN_IN & ~D_REG_14__SCAN_IN & ~D_REG_15__SCAN_IN;
  assign new_n593_ = new_n594_ & new_n595_ & STATE_REG_SCAN_IN & ~new_n270_ & ~new_n534_;
  assign new_n594_ = (IR_REG_22__SCAN_IN | (IR_REG_31__SCAN_IN & (~new_n251_ | ~new_n249_ | ~new_n250_ | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN))) & (~IR_REG_22__SCAN_IN | ~IR_REG_31__SCAN_IN | (new_n251_ & new_n249_ & new_n250_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN)) & (~IR_REG_21__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_20__SCAN_IN & new_n251_ & new_n249_ & new_n250_)));
  assign new_n595_ = (~IR_REG_20__SCAN_IN | IR_REG_31__SCAN_IN) & ((IR_REG_20__SCAN_IN & (~new_n249_ | ~new_n250_ | ~new_n363_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN)) | ~IR_REG_31__SCAN_IN | (~IR_REG_20__SCAN_IN & new_n249_ & new_n250_ & new_n363_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN)) & ((IR_REG_19__SCAN_IN & IR_REG_31__SCAN_IN & (IR_REG_18__SCAN_IN | ~new_n363_ | ~new_n249_ | ~new_n250_)) | (~IR_REG_19__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & new_n249_ & new_n250_ & new_n363_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN));
  assign new_n596_ = (~new_n597_ | (REG3_REG_26__SCAN_IN & new_n393_ & REG3_REG_25__SCAN_IN) | (~REG3_REG_26__SCAN_IN & (~new_n393_ | ~REG3_REG_25__SCAN_IN))) & (~new_n405_ | ~new_n598_) & (STATE_REG_SCAN_IN | ~REG3_REG_26__SCAN_IN);
  assign new_n597_ = STATE_REG_SCAN_IN & ((~new_n584_ & ((new_n252_ ^ ~new_n446_) | (new_n446_ & new_n248_ & ~new_n362_) | (~new_n248_ & ~new_n252_ & new_n446_))) | new_n270_ | new_n534_ | (new_n252_ & ~new_n446_ & (~new_n248_ | new_n362_)));
  assign new_n598_ = new_n599_ & (new_n525_ | (new_n584_ & new_n600_));
  assign new_n599_ = STATE_REG_SCAN_IN & ~new_n270_ & ~new_n534_;
  assign new_n600_ = ~new_n248_ & ~new_n252_ & new_n446_;
  assign new_n601_ = new_n584_ & new_n599_ & ((new_n252_ ^ ~new_n446_) | (new_n446_ & new_n248_ & ~new_n362_));
  assign new_n602_ = new_n649_ & (~new_n603_ | ((new_n488_ | new_n642_ | (~new_n646_ & new_n615_)) & new_n652_ & (~new_n488_ | (~new_n642_ & (new_n646_ | ~new_n615_)))));
  assign new_n603_ = ((~new_n488_ & ~new_n604_ & ~new_n642_) | new_n643_ | (new_n488_ & (new_n604_ | new_n642_))) & (new_n407_ | ~new_n644_) & (~new_n645_ | (new_n616_ & ~new_n488_) | (~new_n616_ & new_n488_));
  assign new_n604_ = new_n615_ & (~new_n612_ | (new_n611_ & (new_n605_ | new_n472_)));
  assign new_n605_ = ~new_n463_ & (~new_n348_ | new_n350_) & ((~new_n348_ & new_n350_) | new_n610_ | (new_n511_ & (new_n318_ | ~new_n322_) & (~new_n606_ | (new_n318_ & ~new_n322_))));
  assign new_n606_ = new_n609_ & (~new_n608_ | (~new_n607_ & (~new_n502_ | (new_n508_ & (~new_n507_ | new_n504_ | new_n506_)))));
  assign new_n607_ = (~new_n306_ | ~new_n310_) & ((new_n287_ & ~new_n291_) | (~new_n306_ & ~new_n310_));
  assign new_n608_ = (~new_n299_ | new_n303_) & (~new_n301_ | new_n307_) & (~new_n327_ | new_n329_) & (~new_n320_ | ~new_n325_);
  assign new_n609_ = (new_n320_ | new_n325_) & ((new_n327_ & ~new_n329_) | (new_n320_ & new_n325_) | ((new_n299_ | ~new_n303_) & (new_n327_ | ~new_n329_) & ((new_n299_ & ~new_n303_) | new_n301_ | ~new_n307_)));
  assign new_n610_ = (~new_n344_ | new_n345_) & ((~new_n339_ & new_n341_) | (~new_n344_ & new_n345_) | (~new_n335_ & new_n336_ & (~new_n339_ | new_n341_)));
  assign new_n611_ = ~new_n516_ & new_n454_ & new_n484_;
  assign new_n612_ = (new_n399_ | new_n401_) & ((new_n399_ & new_n401_) | (~new_n469_ & (~new_n613_ | new_n423_)));
  assign new_n613_ = ~new_n425_ & ((~new_n614_ & ~new_n455_ & ~new_n456_) | new_n487_ | new_n424_ | (new_n426_ & ~new_n455_));
  assign new_n614_ = ((~new_n358_ & DATAI_20_) | (~new_n354_ & new_n356_)) & (new_n360_ | ~new_n361_ | (~new_n358_ & DATAI_20_ & ~new_n354_ & new_n356_));
  assign new_n615_ = ~new_n432_ & (~new_n407_ | ~new_n409_);
  assign new_n616_ = (~new_n407_ | new_n409_) & ((~new_n407_ & new_n409_) | ~new_n641_ | (new_n637_ & ~new_n640_ & ~new_n638_ & (new_n617_ | ~new_n639_)));
  assign new_n617_ = ~new_n632_ & (~new_n630_ | (new_n627_ & (new_n633_ | (new_n636_ & (new_n634_ | new_n618_ | new_n635_)))));
  assign new_n618_ = new_n626_ & (~new_n625_ | (new_n624_ & (~new_n623_ | (~new_n619_ & (~new_n622_ | (new_n620_ & new_n621_))))));
  assign new_n619_ = new_n289_ & ~new_n293_;
  assign new_n620_ = (~new_n272_ | ~new_n277_) & ((~new_n275_ & ~new_n276_) | (~new_n272_ & ~new_n277_));
  assign new_n621_ = ((~new_n261_ & (~new_n283_ | ~new_n284_)) | (~new_n253_ & (~new_n283_ | ~new_n284_))) & (~new_n260_ | ~new_n268_) & (~new_n267_ | new_n273_);
  assign new_n622_ = (((new_n261_ | (new_n283_ & new_n284_)) & (new_n253_ | (new_n283_ & new_n284_))) | ((new_n260_ | new_n268_) & ((new_n260_ & new_n268_) | new_n267_ | ~new_n273_))) & (new_n283_ | new_n284_) & (new_n253_ | new_n261_ | (new_n283_ & new_n284_));
  assign new_n623_ = (new_n287_ | new_n291_) & (new_n289_ | ~new_n293_);
  assign new_n624_ = (~new_n299_ | ~new_n303_) & (~new_n301_ | ~new_n307_) & (~new_n287_ | ~new_n291_) & (~new_n306_ | new_n310_);
  assign new_n625_ = (new_n299_ | new_n303_) & ((new_n299_ & new_n303_) | (new_n301_ & new_n307_) | ((new_n301_ | new_n307_) & (new_n306_ | ~new_n310_)));
  assign new_n626_ = (~new_n327_ | ~new_n329_) & (~new_n318_ | ~new_n322_) & (~new_n320_ | new_n325_);
  assign new_n627_ = (~new_n365_ | new_n368_) & new_n628_ & new_n629_ & (~new_n359_ | ~new_n384_);
  assign new_n628_ = (~new_n360_ | ~new_n361_) & ((~new_n358_ & DATAI_20_) | new_n354_ | ~new_n356_);
  assign new_n629_ = (~new_n344_ | ~new_n345_) & (~new_n348_ | ~new_n350_);
  assign new_n630_ = (new_n365_ | ~new_n368_) & ((new_n365_ & ~new_n368_) | ((new_n353_ | ~new_n357_) & (~new_n628_ | new_n631_)));
  assign new_n631_ = ((new_n359_ & new_n384_) | ((new_n348_ | new_n350_) & (new_n344_ | new_n345_ | (new_n348_ & new_n350_)))) & (new_n359_ | new_n384_) & (new_n360_ | new_n361_);
  assign new_n632_ = new_n370_ & (new_n358_ | ~DATAI_22_);
  assign new_n633_ = ~new_n339_ & ~new_n341_;
  assign new_n634_ = ~new_n335_ & ~new_n336_;
  assign new_n635_ = (~new_n318_ | ~new_n322_) & ((~new_n318_ & ~new_n322_) | (~new_n320_ & new_n325_) | (~new_n327_ & ~new_n329_ & (~new_n318_ | ~new_n322_) & (~new_n320_ | new_n325_)));
  assign new_n636_ = (~new_n335_ | ~new_n336_) & (~new_n339_ | ~new_n341_);
  assign new_n637_ = ~new_n490_ & (~new_n403_ | new_n405_);
  assign new_n638_ = new_n374_ & ~new_n381_;
  assign new_n639_ = (new_n374_ | new_n358_ | ~DATAI_23_) & (new_n370_ | new_n358_ | ~DATAI_22_);
  assign new_n640_ = new_n378_ & ~new_n382_;
  assign new_n641_ = (new_n403_ | ~new_n405_) & (((new_n378_ | ~new_n382_) & (new_n399_ | ~new_n401_)) | (new_n403_ & ~new_n405_) | (new_n399_ & ~new_n401_));
  assign new_n642_ = (~new_n407_ | ~new_n409_) & (new_n421_ | (~new_n407_ & ~new_n409_));
  assign new_n643_ = (new_n248_ | new_n446_) & (~new_n362_ | ~new_n248_ | ~new_n252_);
  assign new_n644_ = new_n594_ & ~new_n262_;
  assign new_n645_ = ~new_n362_ & (new_n248_ | new_n252_) & (~new_n248_ | (new_n252_ ^ ~new_n446_));
  assign new_n646_ = (new_n399_ | new_n401_) & ((new_n399_ & new_n401_) | (new_n648_ & (~new_n647_ | (~new_n605_ & ~new_n472_))));
  assign new_n647_ = new_n454_ & new_n484_;
  assign new_n648_ = ~new_n469_ & (~new_n613_ | new_n423_);
  assign new_n649_ = new_n599_ & (new_n525_ | (new_n650_ & new_n651_));
  assign new_n650_ = (~new_n585_ | ~new_n587_) & (D_REG_1__SCAN_IN | (new_n587_ & new_n586_ & B_REG_SCAN_IN) | new_n585_ | (~new_n586_ & ~B_REG_SCAN_IN)) & (new_n588_ | (new_n587_ & new_n586_ & B_REG_SCAN_IN) | new_n585_ | (~new_n586_ & ~B_REG_SCAN_IN));
  assign new_n651_ = (~new_n594_ | new_n595_) & ((new_n585_ & new_n586_) | (~D_REG_0__SCAN_IN & (~new_n587_ | ~new_n586_ | ~B_REG_SCAN_IN) & ~new_n585_ & (new_n586_ | B_REG_SCAN_IN)));
  assign new_n652_ = ~new_n248_ & new_n252_ & new_n362_;
  assign new_n653_ = ~new_n655_ & ~new_n674_ & ~new_n654_ & (~new_n683_ | (~new_n242_ & ~new_n494_));
  assign new_n654_ = (new_n579_ | new_n576_ | ((new_n577_ | (~new_n578_ ^ ~new_n536_)) & ((~new_n529_ & new_n573_) | (new_n577_ & (new_n578_ | new_n536_) & (~new_n578_ | ~new_n536_))))) & new_n601_ & ((~new_n579_ & ~new_n576_) | (~new_n577_ & (new_n578_ ^ ~new_n536_)) | ((new_n529_ | ~new_n573_) & (~new_n577_ | (~new_n578_ & ~new_n536_) | (new_n578_ & new_n536_))));
  assign new_n655_ = new_n668_ & (((~new_n658_ | (~new_n424_ & ~new_n455_)) & ~new_n672_ & (new_n658_ | new_n424_ | new_n455_)) | ~new_n659_ | ((~new_n656_ | new_n424_ | new_n455_) & ~new_n673_ & (new_n656_ | (~new_n424_ & ~new_n455_))));
  assign new_n656_ = new_n630_ & (new_n657_ | ~new_n627_);
  assign new_n657_ = ~new_n633_ & (~new_n636_ | (~new_n634_ & ~new_n618_ & ~new_n635_));
  assign new_n658_ = ~new_n426_ & (new_n456_ | (new_n614_ & (~new_n484_ | (~new_n605_ & ~new_n472_))));
  assign new_n659_ = new_n666_ & (((~new_n660_ | DATAI_21_) & ~new_n358_ & DATAI_22_) | ~new_n526_ | (new_n660_ & (new_n358_ | ~DATAI_22_) & (new_n358_ | ~DATAI_21_)));
  assign new_n660_ = new_n665_ & new_n384_ & new_n350_ & new_n664_ & new_n336_ & new_n318_ & new_n661_ & new_n663_;
  assign new_n661_ = new_n287_ & ~new_n293_ & new_n284_ & new_n261_ & new_n268_ & ~new_n273_ & new_n662_;
  assign new_n662_ = (~DATAI_1_ | (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_))) & (~new_n278_ | ~new_n262_ | new_n265_ | (new_n263_ & ~new_n264_)) & (~DATAI_0_ | (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_))) & (~IR_REG_0__SCAN_IN | ~new_n262_ | new_n265_ | (new_n263_ & ~new_n264_));
  assign new_n663_ = new_n303_ & new_n307_ & new_n329_ & ~new_n310_ & ~new_n325_;
  assign new_n664_ = new_n341_ & new_n345_;
  assign new_n665_ = new_n361_ & (new_n358_ | ~DATAI_20_);
  assign new_n666_ = (new_n374_ | ~new_n667_) & (new_n365_ | ~new_n644_) & (~new_n600_ | new_n358_ | ~DATAI_22_);
  assign new_n667_ = new_n594_ & new_n262_;
  assign new_n668_ = new_n671_ & ~new_n669_ & new_n599_ & ~new_n670_ & ((~new_n252_ ^ new_n446_) | (~new_n248_ & new_n446_) | (new_n248_ & ~new_n362_));
  assign new_n669_ = (~new_n585_ | ~new_n587_) & (D_REG_1__SCAN_IN | (new_n587_ & new_n586_ & B_REG_SCAN_IN) | new_n585_ | (~new_n586_ & ~B_REG_SCAN_IN));
  assign new_n670_ = ~new_n588_ & (~new_n587_ | ~new_n586_ | ~B_REG_SCAN_IN) & ~new_n585_ & (new_n586_ | B_REG_SCAN_IN);
  assign new_n671_ = (~new_n585_ | ~new_n586_) & (D_REG_0__SCAN_IN | (new_n587_ & new_n586_ & B_REG_SCAN_IN) | new_n585_ | (~new_n586_ & ~B_REG_SCAN_IN));
  assign new_n672_ = (new_n248_ | new_n446_) & (~new_n252_ | ~new_n362_);
  assign new_n673_ = (new_n362_ | (~new_n248_ & ~new_n252_) | (new_n248_ & (~new_n252_ ^ ~new_n446_))) & (~new_n248_ | new_n252_ | ~new_n362_);
  assign new_n674_ = ((~new_n676_ & (new_n493_ | ~new_n421_) & (~new_n493_ | new_n421_)) | ~new_n652_ | (new_n676_ & (new_n493_ ^ new_n421_))) & ~new_n677_ & new_n678_ & ((new_n675_ & new_n493_) | new_n673_ | (~new_n675_ & ~new_n493_));
  assign new_n675_ = new_n641_ & (~new_n637_ | new_n640_ | new_n638_ | (~new_n617_ & new_n639_));
  assign new_n676_ = new_n489_ & ((~new_n399_ & ~new_n401_) | ((~new_n399_ | ~new_n401_) & (~new_n648_ | (new_n647_ & (new_n605_ | new_n472_)))));
  assign new_n677_ = (~new_n493_ | new_n421_ | new_n432_ | (new_n612_ & (~new_n611_ | (~new_n605_ & ~new_n472_)))) & ~new_n643_ & ((new_n493_ & ~new_n421_) | (~new_n493_ & new_n421_) | (~new_n421_ & ~new_n432_ & (~new_n612_ | (new_n611_ & (new_n605_ | new_n472_)))));
  assign new_n678_ = new_n682_ & ((new_n409_ & (new_n405_ | ~new_n679_ | new_n401_)) | ~new_n526_ | (~new_n409_ & ~new_n405_ & new_n679_ & ~new_n401_));
  assign new_n679_ = new_n681_ & new_n660_ & new_n680_;
  assign new_n680_ = (new_n358_ | ~DATAI_22_) & (new_n358_ | ~DATAI_21_);
  assign new_n681_ = ~new_n381_ & ~new_n382_;
  assign new_n682_ = (new_n392_ | ~new_n667_) & (new_n403_ | ~new_n644_) & new_n668_ & (~new_n409_ | ~new_n600_);
  assign new_n683_ = new_n599_ & new_n684_ & new_n594_ & new_n595_;
  assign new_n684_ = ~new_n685_ & ~new_n262_;
  assign new_n685_ = ~new_n265_ & (~new_n263_ | new_n264_);
  assign new_n686_ = (new_n687_ | ~new_n652_) & ~new_n688_ & ~new_n689_ & ~new_n690_ & new_n693_ & (new_n392_ | ~new_n644_);
  assign new_n687_ = ((~new_n642_ & (new_n646_ | ~new_n615_)) | new_n492_ | (new_n392_ & new_n411_)) & ((~new_n646_ & new_n615_) | new_n642_ | ~new_n492_ | (~new_n392_ & ~new_n411_)) & (new_n492_ ? (~new_n392_ | ~new_n411_) : (new_n392_ | new_n411_));
  assign new_n688_ = (new_n492_ | (new_n392_ & ~new_n411_) | (~new_n616_ & (new_n392_ | ~new_n411_))) & ~new_n673_ & (~new_n492_ | ((~new_n392_ | new_n411_) & (new_n616_ | (~new_n392_ & new_n411_))));
  assign new_n689_ = ~new_n643_ & (((new_n604_ | new_n642_) & ~new_n492_ & (~new_n392_ | ~new_n411_)) | (new_n492_ ? (new_n392_ & new_n411_) : (~new_n392_ & ~new_n411_)) | (~new_n604_ & ~new_n642_ & new_n492_ & (new_n392_ | new_n411_)));
  assign new_n690_ = new_n692_ & new_n248_ & (new_n397_ | ~new_n691_ | new_n405_ | ~new_n679_ | new_n401_) & (~new_n397_ | (new_n691_ & ~new_n405_ & new_n679_ & ~new_n401_));
  assign new_n691_ = ~new_n409_ & ~new_n411_;
  assign new_n692_ = ~new_n252_ & new_n446_;
  assign new_n693_ = new_n694_ & (~new_n397_ | ~new_n600_) & (new_n390_ | ~new_n667_ | (~new_n685_ & B_REG_SCAN_IN));
  assign new_n694_ = ~new_n671_ & ~new_n669_ & new_n599_ & ~new_n670_ & ((~new_n252_ ^ new_n446_) | (~new_n248_ & new_n446_) | (new_n248_ & ~new_n362_));
  assign new_n695_ = new_n868_ & ~new_n696_ & new_n863_ & ~new_n700_ & new_n855_ & new_n849_ & new_n721_ & ~new_n878_;
  assign new_n696_ = new_n694_ & (new_n697_ | ~new_n699_ | ((new_n698_ | (~new_n399_ & new_n401_) | (new_n399_ & ~new_n401_)) & ~new_n673_ & (~new_n698_ | (new_n399_ & new_n401_) | (~new_n399_ & ~new_n401_))));
  assign new_n697_ = (~new_n648_ | (new_n647_ & (new_n605_ | new_n472_)) | (new_n399_ ^ new_n401_)) & ~new_n672_ & ((new_n648_ & (~new_n647_ | (~new_n605_ & ~new_n472_))) | (~new_n399_ ^ new_n401_));
  assign new_n698_ = (new_n378_ | ~new_n382_) & ((new_n378_ & ~new_n382_) | new_n638_ | (~new_n617_ & new_n639_));
  assign new_n699_ = ((~new_n679_ & new_n401_) | ~new_n526_ | (new_n679_ & ~new_n401_)) & (new_n403_ | ~new_n667_) & (~new_n401_ | ~new_n600_) & (new_n378_ | ~new_n644_);
  assign new_n700_ = new_n701_ & ((~new_n715_ & (new_n385_ ^ REG2_REG_18__SCAN_IN)) | ~new_n684_ | new_n714_ | (new_n715_ & (new_n385_ | ~REG2_REG_18__SCAN_IN) & (~new_n385_ | REG2_REG_18__SCAN_IN)));
  assign new_n701_ = ((~new_n702_ & (new_n385_ ^ REG1_REG_18__SCAN_IN)) | ~new_n685_ | new_n714_ | (new_n702_ & (new_n385_ | ~REG1_REG_18__SCAN_IN) & (~new_n385_ | REG1_REG_18__SCAN_IN))) & new_n712_ & (new_n714_ | ~new_n262_ | new_n385_);
  assign new_n702_ = (~new_n351_ | REG1_REG_17__SCAN_IN) & ((~new_n351_ & REG1_REG_17__SCAN_IN) | ((new_n346_ | REG1_REG_16__SCAN_IN) & (new_n703_ | (new_n346_ & REG1_REG_16__SCAN_IN))));
  assign new_n703_ = (REG1_REG_15__SCAN_IN | (~new_n337_ & REG1_REG_14__SCAN_IN) | ((~new_n337_ | REG1_REG_14__SCAN_IN) & (new_n704_ | (~new_n319_ & REG1_REG_13__SCAN_IN)))) & (new_n342_ | (REG1_REG_15__SCAN_IN & ((~new_n337_ & REG1_REG_14__SCAN_IN) | ((~new_n337_ | REG1_REG_14__SCAN_IN) & (new_n704_ | (~new_n319_ & REG1_REG_13__SCAN_IN))))));
  assign new_n704_ = new_n711_ & (~new_n710_ | (((~new_n705_ & (~new_n308_ | REG1_REG_9__SCAN_IN)) | (~new_n304_ & REG1_REG_10__SCAN_IN)) & ~new_n709_ & (~new_n304_ | REG1_REG_10__SCAN_IN)));
  assign new_n705_ = new_n708_ & (((new_n706_ | (~new_n294_ & ~REG1_REG_6__SCAN_IN)) & (~new_n288_ | ~REG1_REG_7__SCAN_IN) & (~new_n294_ | ~REG1_REG_6__SCAN_IN)) | (~new_n288_ & ~REG1_REG_7__SCAN_IN) | (~new_n311_ & ~REG1_REG_8__SCAN_IN));
  assign new_n706_ = (~REG1_REG_5__SCAN_IN | ((new_n266_ | ~REG1_REG_4__SCAN_IN) & ((new_n266_ & ~REG1_REG_4__SCAN_IN) | ((~new_n707_ | ~REG1_REG_3__SCAN_IN) & (new_n269_ | (~new_n707_ & ~REG1_REG_3__SCAN_IN)))))) & (~new_n285_ | (~REG1_REG_5__SCAN_IN & (new_n266_ | ~REG1_REG_4__SCAN_IN) & ((new_n266_ & ~REG1_REG_4__SCAN_IN) | ((~new_n707_ | ~REG1_REG_3__SCAN_IN) & (new_n269_ | (~new_n707_ & ~REG1_REG_3__SCAN_IN))))));
  assign new_n707_ = (REG1_REG_2__SCAN_IN | (IR_REG_31__SCAN_IN ? (~IR_REG_2__SCAN_IN ^ (~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN)) : IR_REG_2__SCAN_IN)) & ((REG1_REG_2__SCAN_IN & (IR_REG_2__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_2__SCAN_IN ^ (~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN)))) | (((IR_REG_0__SCAN_IN & REG1_REG_0__SCAN_IN) | (REG1_REG_1__SCAN_IN & (IR_REG_1__SCAN_IN | (IR_REG_0__SCAN_IN & IR_REG_31__SCAN_IN)) & (~IR_REG_1__SCAN_IN | ~IR_REG_0__SCAN_IN | ~IR_REG_31__SCAN_IN))) & (REG1_REG_1__SCAN_IN | (~IR_REG_1__SCAN_IN ^ (~IR_REG_0__SCAN_IN | ~IR_REG_31__SCAN_IN)))));
  assign new_n708_ = (~REG1_REG_8__SCAN_IN | (~IR_REG_8__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & (IR_REG_8__SCAN_IN ^ (new_n249_ & ~IR_REG_7__SCAN_IN)))) & (~REG1_REG_9__SCAN_IN | ((~IR_REG_9__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (new_n249_ & ~IR_REG_7__SCAN_IN & ~IR_REG_8__SCAN_IN & ~IR_REG_9__SCAN_IN) | (IR_REG_9__SCAN_IN & (IR_REG_8__SCAN_IN | ~new_n249_ | IR_REG_7__SCAN_IN)))));
  assign new_n709_ = ~new_n330_ & ~REG1_REG_11__SCAN_IN;
  assign new_n710_ = (~new_n326_ | ~REG1_REG_12__SCAN_IN) & (~new_n330_ | ~REG1_REG_11__SCAN_IN);
  assign new_n711_ = (~new_n319_ | REG1_REG_13__SCAN_IN) & (new_n326_ | REG1_REG_12__SCAN_IN);
  assign new_n712_ = (~new_n713_ | ~ADDR_REG_18__SCAN_IN) & (STATE_REG_SCAN_IN | ~REG3_REG_18__SCAN_IN);
  assign new_n713_ = STATE_REG_SCAN_IN & (new_n270_ | ~new_n534_) & ((~new_n270_ & new_n534_) | (~new_n270_ & new_n594_) | (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)));
  assign new_n714_ = ((~new_n270_ & new_n534_) | (~new_n270_ & new_n594_) | (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)) | ~STATE_REG_SCAN_IN | new_n270_ | new_n534_) & (~new_n270_ | ~STATE_REG_SCAN_IN | (new_n262_ & ~new_n265_ & (~new_n263_ | new_n264_)));
  assign new_n715_ = (~new_n351_ | REG2_REG_17__SCAN_IN) & ((~new_n351_ & REG2_REG_17__SCAN_IN) | ((new_n346_ | REG2_REG_16__SCAN_IN) & ((new_n346_ & REG2_REG_16__SCAN_IN) | ((new_n342_ | REG2_REG_15__SCAN_IN) & (~new_n716_ | (new_n342_ & REG2_REG_15__SCAN_IN))))));
  assign new_n716_ = (new_n337_ | ~REG2_REG_14__SCAN_IN) & ((new_n337_ & ~REG2_REG_14__SCAN_IN) | ((new_n319_ | ~REG2_REG_13__SCAN_IN) & ((new_n319_ & ~REG2_REG_13__SCAN_IN) | ((~new_n326_ | ~REG2_REG_12__SCAN_IN) & (new_n717_ | (~new_n326_ & ~REG2_REG_12__SCAN_IN))))));
  assign new_n717_ = (~new_n330_ | ~REG2_REG_11__SCAN_IN) & ((~new_n330_ & ~REG2_REG_11__SCAN_IN) | ((new_n304_ | ~REG2_REG_10__SCAN_IN) & ((new_n304_ & ~REG2_REG_10__SCAN_IN) | ((new_n308_ | ~REG2_REG_9__SCAN_IN) & (new_n718_ | (new_n308_ & ~REG2_REG_9__SCAN_IN))))));
  assign new_n718_ = (~new_n311_ | ~REG2_REG_8__SCAN_IN) & ((~new_n311_ & ~REG2_REG_8__SCAN_IN) | ((~new_n288_ | ~REG2_REG_7__SCAN_IN) & ((~new_n719_ & (~new_n294_ | ~REG2_REG_6__SCAN_IN)) | (~new_n288_ & ~REG2_REG_7__SCAN_IN) | (~new_n294_ & ~REG2_REG_6__SCAN_IN))));
  assign new_n719_ = (new_n285_ | REG2_REG_5__SCAN_IN) & ((new_n285_ & REG2_REG_5__SCAN_IN) | (~new_n266_ & REG2_REG_4__SCAN_IN) | ((~new_n266_ | REG2_REG_4__SCAN_IN) & ((~new_n269_ & REG2_REG_3__SCAN_IN) | (~new_n720_ & (~new_n269_ | REG2_REG_3__SCAN_IN)))));
  assign new_n720_ = (~REG2_REG_2__SCAN_IN | (~IR_REG_2__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & (IR_REG_2__SCAN_IN ^ (~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN)))) & ((~REG2_REG_2__SCAN_IN & (IR_REG_31__SCAN_IN ? (IR_REG_2__SCAN_IN ^ (~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN)) : ~IR_REG_2__SCAN_IN)) | ((~IR_REG_0__SCAN_IN | ~REG2_REG_0__SCAN_IN) & (~REG2_REG_1__SCAN_IN | (~IR_REG_1__SCAN_IN & (~IR_REG_0__SCAN_IN | ~IR_REG_31__SCAN_IN)) | (IR_REG_1__SCAN_IN & IR_REG_0__SCAN_IN & IR_REG_31__SCAN_IN))) | (~REG2_REG_1__SCAN_IN & (IR_REG_1__SCAN_IN ^ (~IR_REG_0__SCAN_IN | ~IR_REG_31__SCAN_IN))));
  assign new_n721_ = ~new_n842_ & ~new_n845_ & ~new_n722_ & ~new_n724_ & new_n837_ & ~new_n728_ & new_n733_ & new_n812_;
  assign new_n722_ = (~new_n411_ | (~new_n409_ & ~new_n405_ & new_n679_ & ~new_n401_)) & new_n723_ & (new_n409_ | new_n411_ | new_n405_ | ~new_n679_ | new_n401_);
  assign new_n723_ = new_n692_ & new_n595_ & new_n599_ & (new_n525_ | (new_n650_ & new_n651_));
  assign new_n724_ = new_n668_ & (((new_n725_ | new_n482_) & ~new_n672_ & (~new_n725_ | ~new_n482_)) | ~new_n726_ | ((new_n482_ | (~new_n618_ & ~new_n635_)) & ~new_n673_ & (~new_n482_ | new_n618_ | new_n635_)));
  assign new_n725_ = (new_n318_ | ~new_n322_) & (~new_n606_ | (new_n318_ & ~new_n322_));
  assign new_n726_ = ((~new_n727_ & ~new_n336_) | ~new_n526_ | (new_n727_ & new_n336_)) & (new_n339_ | ~new_n667_) & (new_n336_ | ~new_n600_) & (new_n322_ | ~new_n644_);
  assign new_n727_ = new_n318_ & new_n661_ & new_n663_;
  assign new_n728_ = new_n730_ & ((new_n729_ & ~new_n560_ & ~new_n561_) | ~new_n601_ | (~new_n729_ & (new_n560_ | new_n561_)));
  assign new_n729_ = ~new_n562_ & (new_n531_ | ~new_n547_);
  assign new_n730_ = (new_n731_ | (~new_n302_ & ~REG3_REG_9__SCAN_IN) | (new_n302_ & REG3_REG_9__SCAN_IN)) & ~new_n732_ & (STATE_REG_SCAN_IN | ~REG3_REG_9__SCAN_IN) & (~new_n598_ | new_n307_);
  assign new_n731_ = (~STATE_REG_SCAN_IN | ((new_n584_ | ((~new_n252_ ^ ~new_n446_) & (~new_n446_ | ~new_n248_ | new_n362_) & (new_n248_ | new_n252_ | ~new_n446_))) & ~new_n270_ & ~new_n534_ & (~new_n252_ | new_n446_ | (new_n248_ & ~new_n362_)))) & (new_n584_ | ~STATE_REG_SCAN_IN | new_n270_ | new_n534_ | ~new_n252_ | new_n446_ | ~new_n248_ | new_n362_);
  assign new_n732_ = new_n593_ & ((~new_n306_ & new_n584_ & ~new_n262_) | (~new_n299_ & new_n584_ & new_n262_));
  assign new_n733_ = new_n805_ & ~new_n734_ & ~new_n738_ & ~new_n811_ & new_n744_ & new_n798_;
  assign new_n734_ = new_n649_ & (((~new_n736_ | new_n737_) & ~new_n672_ & (new_n736_ | ~new_n737_)) | (~new_n283_ & new_n644_) | (new_n645_ & (new_n735_ | ~new_n737_) & (~new_n735_ | new_n737_)));
  assign new_n735_ = new_n622_ & (~new_n620_ | ~new_n621_);
  assign new_n736_ = (~new_n283_ | new_n284_) & ((~new_n506_ & (~new_n253_ | new_n261_)) | (~new_n253_ & new_n261_) | (~new_n283_ & new_n284_));
  assign new_n737_ = ~new_n289_ ^ new_n293_;
  assign new_n738_ = new_n739_ & ((~new_n743_ & ~new_n742_ & (new_n741_ | new_n539_ | (~new_n540_ & ~new_n541_))) | ~new_n601_ | (new_n743_ & (new_n742_ | (~new_n741_ & ~new_n539_ & (new_n540_ | new_n541_)))));
  assign new_n739_ = (new_n731_ | REG3_REG_3__SCAN_IN) & new_n740_ & (~new_n593_ | ((new_n253_ | ~new_n584_ | ~new_n262_) & (new_n267_ | ~new_n584_ | new_n262_)));
  assign new_n740_ = (STATE_REG_SCAN_IN | ~REG3_REG_3__SCAN_IN) & (new_n268_ | ~new_n599_ | (~new_n525_ & (~new_n584_ | ~new_n600_)));
  assign new_n741_ = (new_n536_ | ((new_n267_ | ~new_n533_) & (~new_n273_ | ~new_n535_))) & (~new_n536_ | (~new_n267_ & new_n533_) | (new_n273_ & new_n535_)) & (new_n267_ | ~new_n537_) & (~new_n273_ | ~new_n533_);
  assign new_n742_ = (new_n536_ ^ ((~new_n267_ & new_n533_) | (new_n273_ & new_n535_))) & ((~new_n267_ & new_n537_) | (new_n273_ & new_n533_));
  assign new_n743_ = ((~new_n260_ & new_n537_) | (~new_n268_ & new_n533_)) ^ (new_n536_ ^ ((~new_n260_ & new_n533_) | (~new_n268_ & new_n535_)));
  assign new_n744_ = new_n783_ & new_n745_ & new_n782_ & new_n756_ & new_n761_ & ~new_n790_ & ~new_n791_ & new_n793_;
  assign new_n745_ = (~new_n597_ | ~new_n259_) & (~new_n598_ | new_n746_) & ~new_n747_ & (~new_n754_ | new_n755_);
  assign new_n746_ = new_n261_ & ~new_n381_ & ~new_n273_ & new_n303_;
  assign new_n747_ = (new_n714_ | (~new_n748_ & ~new_n750_ & ~new_n751_)) & (STATE_REG_SCAN_IN | ~REG3_REG_5__SCAN_IN) & (~new_n713_ | ~ADDR_REG_5__SCAN_IN);
  assign new_n748_ = (~new_n749_ | ~new_n285_) & (new_n749_ | new_n285_) & ~new_n265_ & (~new_n263_ | new_n264_);
  assign new_n749_ = REG1_REG_5__SCAN_IN ^ ((~new_n266_ & REG1_REG_4__SCAN_IN) | ((~new_n266_ | REG1_REG_4__SCAN_IN) & ((new_n707_ & REG1_REG_3__SCAN_IN) | (~new_n269_ & (new_n707_ | REG1_REG_3__SCAN_IN)))));
  assign new_n750_ = new_n262_ & new_n285_;
  assign new_n751_ = ~new_n752_ & ~new_n753_ & ~new_n262_ & (new_n265_ | (new_n263_ & ~new_n264_));
  assign new_n752_ = (~new_n285_ | ~REG2_REG_5__SCAN_IN) & (new_n285_ | REG2_REG_5__SCAN_IN) & ((~new_n266_ & REG2_REG_4__SCAN_IN) | ((~new_n266_ | REG2_REG_4__SCAN_IN) & ((~new_n269_ & REG2_REG_3__SCAN_IN) | (~new_n720_ & (~new_n269_ | REG2_REG_3__SCAN_IN)))));
  assign new_n753_ = (~new_n285_ ^ REG2_REG_5__SCAN_IN) & (new_n266_ | ~REG2_REG_4__SCAN_IN) & ((new_n266_ & ~REG2_REG_4__SCAN_IN) | ((new_n269_ | ~REG2_REG_3__SCAN_IN) & (new_n720_ | (new_n269_ & ~REG2_REG_3__SCAN_IN))));
  assign new_n754_ = new_n667_ & new_n599_ & (new_n525_ | (new_n650_ & new_n651_));
  assign new_n755_ = new_n360_ & new_n291_ & new_n335_;
  assign new_n756_ = (new_n668_ | new_n758_) & (new_n694_ | new_n760_) & (~new_n668_ | new_n757_) & (new_n668_ | ~REG1_REG_0__SCAN_IN);
  assign new_n757_ = ((new_n672_ & new_n673_) | (~new_n275_ ^ new_n276_)) & (new_n275_ | ~new_n692_) & (new_n272_ | ~new_n667_);
  assign new_n758_ = new_n759_ & REG1_REG_30__SCAN_IN & REG1_REG_26__SCAN_IN & REG1_REG_27__SCAN_IN;
  assign new_n759_ = ~REG1_REG_3__SCAN_IN & REG1_REG_4__SCAN_IN & REG1_REG_13__SCAN_IN & ~REG1_REG_14__SCAN_IN & REG1_REG_17__SCAN_IN & ~REG1_REG_22__SCAN_IN;
  assign new_n760_ = ~REG0_REG_1__SCAN_IN & ~REG0_REG_7__SCAN_IN & ~REG0_REG_24__SCAN_IN & ~REG0_REG_25__SCAN_IN & REG0_REG_29__SCAN_IN & ~REG0_REG_31__SCAN_IN;
  assign new_n761_ = ~new_n762_ & ~new_n765_ & (~new_n763_ | (new_n344_ & ~new_n299_ & new_n320_)) & new_n767_ & (~new_n359_ | ~new_n763_);
  assign new_n762_ = (new_n763_ | ~new_n764_) & (~new_n253_ | ~new_n291_ | ~new_n763_ | new_n301_ | ~new_n327_);
  assign new_n763_ = STATE_REG_SCAN_IN & ~new_n270_ & new_n534_;
  assign new_n764_ = ~DATAO_REG_7__SCAN_IN & DATAO_REG_9__SCAN_IN & DATAO_REG_20__SCAN_IN & DATAO_REG_10__SCAN_IN & ~DATAO_REG_16__SCAN_IN;
  assign new_n765_ = (new_n714_ | new_n766_) & (STATE_REG_SCAN_IN | ~REG3_REG_0__SCAN_IN) & (~new_n713_ | ~ADDR_REG_0__SCAN_IN);
  assign new_n766_ = ((~IR_REG_0__SCAN_IN & ~REG2_REG_0__SCAN_IN) | (IR_REG_0__SCAN_IN & REG2_REG_0__SCAN_IN) | new_n262_ | (~new_n265_ & (~new_n263_ | new_n264_))) & (~new_n262_ | ~IR_REG_0__SCAN_IN) & (new_n265_ | (new_n263_ & ~new_n264_) | (~IR_REG_0__SCAN_IN & ~REG1_REG_0__SCAN_IN) | (IR_REG_0__SCAN_IN & REG1_REG_0__SCAN_IN));
  assign new_n767_ = ~new_n769_ & new_n781_ & ~new_n772_ & new_n773_ & (~B_REG_SCAN_IN | (new_n768_ & new_n771_));
  assign new_n768_ = STATE_REG_SCAN_IN & (new_n270_ | ~new_n534_);
  assign new_n769_ = new_n362_ & new_n526_ & STATE_REG_SCAN_IN & ~new_n270_ & ~new_n534_ & (~new_n770_ | (new_n355_ ^ REG3_REG_18__SCAN_IN));
  assign new_n770_ = ~new_n290_ & (~REG3_REG_13__SCAN_IN ^ (REG3_REG_12__SCAN_IN & new_n321_ & REG3_REG_11__SCAN_IN));
  assign new_n771_ = new_n270_ ? ~new_n252_ : (new_n595_ & new_n252_ & ~new_n446_ & ~new_n262_ & (new_n265_ | (new_n263_ & ~new_n264_)));
  assign new_n772_ = ((new_n587_ & new_n586_ & B_REG_SCAN_IN) | new_n585_ | (~new_n586_ & ~B_REG_SCAN_IN)) & STATE_REG_SCAN_IN & ~new_n270_ & ~new_n534_;
  assign new_n773_ = ~new_n776_ & new_n777_ & ((~new_n774_ & new_n775_) | ~STATE_REG_SCAN_IN | ~IR_REG_31__SCAN_IN);
  assign new_n774_ = ~IR_REG_12__SCAN_IN ^ (~IR_REG_11__SCAN_IN & ~IR_REG_10__SCAN_IN & new_n305_ & new_n249_ & ~IR_REG_7__SCAN_IN);
  assign new_n775_ = ((IR_REG_16__SCAN_IN & (IR_REG_15__SCAN_IN | IR_REG_14__SCAN_IN | ~new_n249_ | ~new_n250_)) | (~IR_REG_15__SCAN_IN & ~IR_REG_16__SCAN_IN & ~IR_REG_14__SCAN_IN & new_n249_ & new_n250_)) & (new_n249_ | new_n295_) & (~IR_REG_8__SCAN_IN ^ (~new_n249_ | IR_REG_7__SCAN_IN));
  assign new_n776_ = (~STATE_REG_SCAN_IN | ~IR_REG_31__SCAN_IN | (~IR_REG_15__SCAN_IN & ~IR_REG_14__SCAN_IN & new_n249_ & new_n250_) | (IR_REG_15__SCAN_IN & (IR_REG_14__SCAN_IN | ~new_n249_ | ~new_n250_))) & (~DATAI_15_ | STATE_REG_SCAN_IN) & (IR_REG_31__SCAN_IN | ~STATE_REG_SCAN_IN | ~IR_REG_15__SCAN_IN);
  assign new_n777_ = new_n780_ & ((~new_n778_ & STATE_REG_SCAN_IN) | (new_n779_ & ~REG3_REG_23__SCAN_IN & ~REG3_REG_10__SCAN_IN & ~REG3_REG_4__SCAN_IN & ~REG3_REG_2__SCAN_IN));
  assign new_n778_ = (~IR_REG_31__SCAN_IN | (~IR_REG_2__SCAN_IN ^ (~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN))) & (IR_REG_2__SCAN_IN | IR_REG_31__SCAN_IN | IR_REG_6__SCAN_IN | IR_REG_8__SCAN_IN | IR_REG_12__SCAN_IN | IR_REG_16__SCAN_IN);
  assign new_n779_ = ~DATAI_16_ & ~DATAI_12_ & ~DATAI_2_ & ~STATE_REG_SCAN_IN & ~DATAI_8_ & ~DATAI_6_;
  assign new_n780_ = ~D_REG_22__SCAN_IN & D_REG_27__SCAN_IN & D_REG_11__SCAN_IN & ~D_REG_19__SCAN_IN;
  assign new_n781_ = ((STATE_REG_SCAN_IN & ~new_n270_ & new_n534_) | (~DATAO_REG_12__SCAN_IN & ~DATAO_REG_4__SCAN_IN & ~DATAO_REG_11__SCAN_IN)) & (DATAO_REG_18__SCAN_IN | (STATE_REG_SCAN_IN & ~new_n270_ & new_n534_));
  assign new_n782_ = (~new_n353_ | ~new_n763_) & (~new_n649_ | ~new_n600_ | (new_n384_ & ~new_n293_ & ~new_n411_));
  assign new_n783_ = ~new_n786_ & (~new_n784_ | (new_n737_ & (~new_n622_ | (new_n620_ & new_n621_))) | (~new_n737_ & new_n622_ & (~new_n620_ | ~new_n621_)));
  assign new_n784_ = new_n785_ & new_n599_ & (new_n525_ | (new_n650_ & new_n651_));
  assign new_n785_ = new_n248_ & ~new_n446_ & new_n362_;
  assign new_n786_ = ~new_n788_ & STATE_REG_SCAN_IN & (~new_n787_ | (~new_n584_ & ((~new_n252_ ^ new_n446_) | (new_n446_ & new_n248_ & ~new_n362_) | (~new_n248_ & ~new_n252_ & new_n446_))));
  assign new_n787_ = ~new_n270_ & ~new_n534_ & (~new_n594_ | new_n595_);
  assign new_n788_ = new_n789_ & (~REG3_REG_23__SCAN_IN ^ (REG3_REG_22__SCAN_IN & REG3_REG_21__SCAN_IN & REG3_REG_20__SCAN_IN & REG3_REG_19__SCAN_IN & new_n355_ & REG3_REG_18__SCAN_IN));
  assign new_n789_ = ~REG3_REG_2__SCAN_IN & (new_n300_ ^ ~REG3_REG_10__SCAN_IN);
  assign new_n790_ = new_n601_ & ((~new_n741_ & ~new_n742_) ^ (~new_n539_ & (new_n540_ | new_n541_)));
  assign new_n791_ = new_n694_ & ((((~new_n275_ & new_n276_) | (~new_n272_ & new_n277_) | (new_n272_ & ~new_n277_)) & ~new_n672_ & (new_n275_ | ~new_n276_ | (~new_n272_ ^ new_n277_))) | ~new_n792_ | ((new_n275_ | new_n276_ | (~new_n272_ ^ new_n277_)) & ~new_n673_ & ((~new_n275_ & ~new_n276_) | (~new_n272_ & new_n277_) | (new_n272_ & ~new_n277_))));
  assign new_n792_ = ((~new_n275_ & ~new_n277_) | ~new_n526_ | (new_n275_ & new_n277_)) & (new_n267_ | ~new_n667_) & (new_n277_ | ~new_n600_) & (new_n276_ | ~new_n644_);
  assign new_n793_ = ~new_n795_ & ~new_n796_ & ~new_n797_ & ((~new_n794_ & new_n293_) | ~new_n723_ | (new_n794_ & ~new_n293_));
  assign new_n794_ = new_n284_ & new_n261_ & new_n268_ & ~new_n273_ & new_n662_;
  assign new_n795_ = (REG2_REG_6__SCAN_IN | REG2_REG_13__SCAN_IN | REG2_REG_18__SCAN_IN | REG2_REG_28__SCAN_IN) & (~new_n599_ | (~new_n525_ & (~new_n650_ | ~new_n651_)));
  assign new_n796_ = (~new_n584_ | ((~new_n327_ | ~new_n260_ | ~new_n262_) & (~new_n301_ | ~new_n272_ | new_n262_))) & new_n593_ & (new_n584_ | ~new_n789_);
  assign new_n797_ = ~new_n318_ & new_n600_ & new_n599_ & (new_n525_ | (new_n650_ & new_n651_));
  assign new_n798_ = (~new_n801_ | (new_n649_ & (~new_n799_ | new_n804_))) & (~new_n723_ | (new_n318_ & new_n661_ & new_n663_) | (~new_n318_ & (~new_n661_ | ~new_n663_)));
  assign new_n799_ = (new_n800_ | ~new_n645_) & (new_n272_ | ~new_n644_);
  assign new_n800_ = ((new_n272_ & new_n277_) | ((new_n275_ | new_n276_) & (new_n272_ | new_n277_))) ^ (~new_n267_ ^ new_n273_);
  assign new_n801_ = new_n802_ & (~new_n784_ | new_n800_) & (~new_n754_ | new_n260_) & (~new_n723_ | (new_n273_ & ~new_n662_) | (~new_n273_ & new_n662_));
  assign new_n802_ = (~new_n273_ | ~new_n600_ | ~new_n599_ | (~new_n525_ & (~new_n650_ | ~new_n651_))) & ~new_n803_ & (~REG2_REG_2__SCAN_IN | (new_n599_ & (new_n525_ | (new_n650_ & new_n651_))));
  assign new_n803_ = REG3_REG_2__SCAN_IN & new_n362_ & new_n526_ & STATE_REG_SCAN_IN & ~new_n270_ & ~new_n534_;
  assign new_n804_ = ((new_n272_ & ~new_n277_) | (~new_n275_ & new_n276_ & (new_n272_ | ~new_n277_)) | (~new_n267_ ^ new_n273_)) & ~new_n672_ & (((~new_n272_ | new_n277_) & (new_n275_ | ~new_n276_ | (~new_n272_ & new_n277_))) | (~new_n267_ & new_n273_) | (new_n267_ & ~new_n273_));
  assign new_n805_ = ((~new_n806_ & ~new_n384_) | ~new_n723_ | (new_n806_ & new_n384_)) & (~new_n694_ | (~new_n807_ & ~new_n808_ & new_n809_));
  assign new_n806_ = new_n350_ & new_n664_ & new_n336_ & new_n318_ & new_n661_ & new_n663_;
  assign new_n807_ = ((~new_n287_ & ~new_n291_) | (new_n287_ & new_n291_) | ~new_n508_ | (new_n507_ & ~new_n504_ & ~new_n506_)) & ~new_n672_ & ((~new_n287_ ^ ~new_n291_) | (new_n508_ & (~new_n507_ | new_n504_ | new_n506_)));
  assign new_n808_ = ((new_n287_ ^ new_n291_) | (~new_n289_ & new_n293_) | ((~new_n289_ | new_n293_) & (~new_n622_ | (new_n620_ & new_n621_)))) & ~new_n673_ & ((new_n287_ & new_n291_) | (~new_n287_ & ~new_n291_) | ((new_n289_ | ~new_n293_) & ((new_n289_ & ~new_n293_) | (new_n622_ & (~new_n620_ | ~new_n621_)))));
  assign new_n809_ = ((~new_n810_ & ~new_n287_) | ~new_n692_ | ~new_n248_ | (new_n810_ & new_n287_)) & (new_n306_ | ~new_n667_) & (new_n289_ | ~new_n644_) & (new_n287_ | ~new_n692_ | new_n248_);
  assign new_n810_ = ~new_n293_ & new_n284_ & new_n261_ & new_n268_ & ~new_n273_ & new_n662_;
  assign new_n811_ = new_n525_ & new_n599_ & (REG3_REG_28__SCAN_IN | (REG3_REG_27__SCAN_IN & REG3_REG_26__SCAN_IN & new_n393_ & REG3_REG_25__SCAN_IN)) & (~REG3_REG_28__SCAN_IN | ~REG3_REG_27__SCAN_IN | ~REG3_REG_26__SCAN_IN | ~new_n393_ | ~REG3_REG_25__SCAN_IN);
  assign new_n812_ = ~new_n813_ & ~new_n818_ & new_n825_ & ~new_n823_ & (new_n395_ | ~new_n754_);
  assign new_n813_ = new_n784_ & (~new_n477_ ^ (~new_n816_ & (new_n814_ | ~new_n817_)));
  assign new_n814_ = ~new_n815_ & (~new_n625_ | (new_n624_ & (~new_n623_ | (~new_n619_ & (~new_n622_ | (new_n620_ & new_n621_))))));
  assign new_n815_ = new_n327_ & new_n329_;
  assign new_n816_ = new_n320_ & ~new_n325_;
  assign new_n817_ = (new_n320_ | ~new_n325_) & (new_n327_ | new_n329_);
  assign new_n818_ = new_n820_ & (~new_n601_ | (~new_n822_ ^ (new_n548_ | (new_n546_ & (~new_n819_ | new_n538_)))));
  assign new_n819_ = ~new_n545_ & (~new_n544_ | new_n539_ | (~new_n540_ & ~new_n541_));
  assign new_n820_ = (new_n731_ | ~new_n290_) & new_n821_ & (~new_n593_ | ((new_n291_ | ~new_n584_ | ~new_n262_) & (new_n283_ | ~new_n584_ | new_n262_)));
  assign new_n821_ = (STATE_REG_SCAN_IN | ~REG3_REG_6__SCAN_IN) & (~new_n293_ | ~new_n599_ | (~new_n525_ & (~new_n584_ | ~new_n600_)));
  assign new_n822_ = (~new_n536_ ^ ((~new_n289_ & new_n533_) | (new_n293_ & new_n535_))) ^ ((new_n289_ | ~new_n537_) & (~new_n293_ | ~new_n533_));
  assign new_n823_ = (new_n824_ | ~new_n584_) & new_n593_ & (new_n375_ | new_n584_ | new_n259_);
  assign new_n824_ = (~new_n370_ | ~new_n260_ | new_n262_) & (~new_n378_ | ~new_n283_ | ~new_n262_);
  assign new_n825_ = ((~new_n835_ & (~new_n819_ | ~new_n836_) & (new_n819_ | new_n836_)) | ~new_n601_ | (new_n835_ & (~new_n819_ ^ new_n836_))) & (~new_n668_ | (~new_n826_ & new_n830_));
  assign new_n826_ = ((new_n506_ & (new_n253_ ^ new_n261_)) | new_n672_ | (~new_n506_ & (new_n253_ | ~new_n261_) & (~new_n253_ | new_n261_))) & ~new_n828_ & new_n829_ & ((new_n827_ & (new_n253_ | ~new_n261_) & (~new_n253_ | new_n261_)) | new_n673_ | (~new_n827_ & (new_n253_ ^ new_n261_)));
  assign new_n827_ = (new_n260_ | new_n268_) & ((new_n260_ & new_n268_) | ((new_n267_ | ~new_n273_) & ((new_n272_ & new_n277_) | ((new_n275_ | new_n276_) & (new_n272_ | new_n277_)) | (new_n267_ & ~new_n273_))));
  assign new_n828_ = (new_n261_ | (new_n268_ & ~new_n273_ & new_n662_)) & new_n526_ & (~new_n261_ | ~new_n268_ | new_n273_ | ~new_n662_);
  assign new_n829_ = (new_n283_ | ~new_n667_) & (new_n260_ | ~new_n644_) & (new_n261_ | ~new_n600_);
  assign new_n830_ = ((new_n832_ & (~new_n260_ | new_n268_) & (new_n260_ | ~new_n268_)) | new_n673_ | (~new_n832_ & (~new_n260_ ^ ~new_n268_))) & new_n833_ & ((new_n831_ & (~new_n260_ | new_n268_) & (new_n260_ | ~new_n268_)) | new_n672_ | (~new_n831_ & (~new_n260_ ^ ~new_n268_)));
  assign new_n831_ = (~new_n267_ | ~new_n273_) & ((~new_n267_ & ~new_n273_) | ((~new_n272_ | new_n277_) & (new_n275_ | ~new_n276_ | (~new_n272_ & new_n277_))));
  assign new_n832_ = (new_n267_ | ~new_n273_) & ((new_n267_ & ~new_n273_) | (new_n272_ & new_n277_) | ((new_n275_ | new_n276_) & (new_n272_ | new_n277_)));
  assign new_n833_ = ((~new_n268_ & (new_n273_ | ~new_n662_)) | ~new_n526_ | (new_n268_ & ~new_n273_ & new_n662_)) & ~new_n834_ & (new_n267_ | ~new_n644_) & (new_n268_ | ~new_n600_);
  assign new_n834_ = new_n594_ & new_n262_ & ((REG1_REG_4__SCAN_IN & ~new_n254_ & ~new_n257_) | (REG0_REG_4__SCAN_IN & new_n254_ & ~new_n257_) | (new_n259_ & ~new_n254_ & new_n257_) | (REG2_REG_4__SCAN_IN & new_n254_ & new_n257_));
  assign new_n835_ = (new_n253_ | ~new_n537_) & (new_n261_ | ~new_n533_);
  assign new_n836_ = ~new_n536_ ^ ((~new_n253_ & new_n533_) | (~new_n261_ & new_n535_));
  assign new_n837_ = (~new_n838_ | ~new_n840_) & ((~new_n554_ & ~new_n556_ & ~new_n560_ & (new_n729_ | new_n561_)) | ~new_n601_ | ((new_n554_ | new_n556_) & (new_n560_ | (~new_n729_ & ~new_n561_))));
  assign new_n838_ = ((new_n606_ & ~new_n477_) | new_n672_ | (~new_n606_ & new_n477_)) & ~new_n839_ & (~new_n645_ | (new_n477_ ^ (~new_n816_ & (new_n814_ | ~new_n817_))));
  assign new_n839_ = ~new_n320_ & new_n644_;
  assign new_n840_ = new_n841_ & (~new_n248_ | new_n252_ | ~new_n362_ | (new_n477_ ^ (~new_n816_ & (new_n814_ | ~new_n817_))));
  assign new_n841_ = (~new_n526_ | (new_n318_ & new_n661_ & new_n663_) | (~new_n318_ & (~new_n661_ | ~new_n663_))) & new_n668_ & (new_n318_ | ~new_n600_) & (new_n335_ | ~new_n667_);
  assign new_n842_ = new_n649_ & (~new_n838_ | (new_n785_ & (~new_n844_ ^ (~new_n843_ | (~new_n657_ & new_n629_)))));
  assign new_n843_ = (new_n348_ | new_n350_) & (new_n344_ | new_n345_ | (new_n348_ & new_n350_));
  assign new_n844_ = ~new_n359_ ^ new_n384_;
  assign new_n845_ = ~new_n846_ & new_n847_ & (((new_n348_ | ~new_n350_) & (~new_n348_ | new_n350_) & (new_n344_ | new_n345_) & (new_n657_ | (new_n344_ & new_n345_))) | new_n673_ | ((new_n348_ ^ new_n350_) & ((~new_n344_ & ~new_n345_) | (~new_n657_ & (~new_n344_ | ~new_n345_)))));
  assign new_n846_ = ((~new_n348_ ^ new_n350_) | new_n610_ | (new_n511_ & (new_n318_ | ~new_n322_) & (~new_n606_ | (new_n318_ & ~new_n322_)))) & ~new_n672_ & ((~new_n348_ & new_n350_) | (new_n348_ & ~new_n350_) | (~new_n610_ & (~new_n511_ | (~new_n318_ & new_n322_) | (new_n606_ & (~new_n318_ | new_n322_)))));
  assign new_n847_ = ~new_n848_ & (new_n359_ | ~new_n667_) & new_n668_ & (new_n350_ | ~new_n600_) & (new_n344_ | ~new_n644_);
  assign new_n848_ = (new_n350_ | (new_n664_ & new_n336_ & new_n318_ & new_n661_ & new_n663_)) & new_n526_ & (~new_n350_ | ~new_n664_ | ~new_n336_ | ~new_n318_ | ~new_n661_ | ~new_n663_);
  assign new_n849_ = ((~new_n389_ & new_n850_ & new_n692_) | ~new_n668_ | new_n854_ | (~new_n850_ & new_n389_ & new_n692_)) & (~new_n852_ | (~new_n851_ & new_n601_));
  assign new_n850_ = new_n248_ & (new_n397_ | ~new_n691_ | new_n405_ | ~new_n679_ | new_n401_);
  assign new_n851_ = (~new_n530_ & ~new_n570_) ^ (~new_n569_ & ~new_n571_);
  assign new_n852_ = (new_n731_ | (~new_n340_ & ~REG3_REG_15__SCAN_IN) | (new_n340_ & REG3_REG_15__SCAN_IN)) & ~new_n853_ & (STATE_REG_SCAN_IN | ~REG3_REG_15__SCAN_IN) & (~new_n598_ | new_n341_);
  assign new_n853_ = new_n593_ & ((~new_n335_ & new_n584_ & ~new_n262_) | (~new_n344_ & new_n584_ & new_n262_));
  assign new_n854_ = ~new_n391_ & new_n667_ & (new_n685_ | ~B_REG_SCAN_IN);
  assign new_n855_ = ~new_n857_ & ~new_n861_ & (~new_n649_ | (new_n860_ & ((~new_n856_ & ~new_n844_) | new_n672_ | (new_n856_ & new_n844_))));
  assign new_n856_ = (~new_n348_ | new_n350_) & ((~new_n348_ & new_n350_) | new_n610_ | (new_n725_ & new_n511_));
  assign new_n857_ = (new_n714_ | (~new_n858_ & new_n859_)) & (~new_n713_ | ~ADDR_REG_16__SCAN_IN) & (STATE_REG_SCAN_IN | ~REG3_REG_16__SCAN_IN);
  assign new_n858_ = ((new_n346_ & REG2_REG_16__SCAN_IN) | (~new_n346_ & ~REG2_REG_16__SCAN_IN) | (~new_n342_ & ~REG2_REG_15__SCAN_IN) | (new_n716_ & (~new_n342_ | ~REG2_REG_15__SCAN_IN))) & new_n684_ & ((new_n346_ ^ REG2_REG_16__SCAN_IN) | ((new_n342_ | REG2_REG_15__SCAN_IN) & (~new_n716_ | (new_n342_ & REG2_REG_15__SCAN_IN))));
  assign new_n859_ = (~new_n262_ | ~new_n346_) & ((new_n703_ & (new_n346_ | REG1_REG_16__SCAN_IN) & (~new_n346_ | ~REG1_REG_16__SCAN_IN)) | ~new_n685_ | (~new_n703_ & (new_n346_ ^ ~REG1_REG_16__SCAN_IN)));
  assign new_n860_ = (new_n348_ | ~new_n644_) & (~new_n645_ | (new_n844_ ^ (~new_n843_ | (~new_n657_ & new_n629_))));
  assign new_n861_ = new_n694_ & (((~new_n862_ | (~new_n358_ & DATAI_31_)) & new_n526_ & (new_n862_ | new_n358_ | ~DATAI_31_)) | new_n854_ | (new_n600_ & ~new_n358_ & DATAI_31_));
  assign new_n862_ = ~new_n389_ & ~new_n397_ & new_n691_ & ~new_n405_ & ~new_n401_ & new_n681_ & new_n660_ & new_n680_;
  assign new_n863_ = (new_n864_ | ~new_n866_) & (~new_n784_ | (~new_n616_ & new_n488_) | (new_n616_ & ~new_n488_));
  assign new_n864_ = new_n601_ & (new_n865_ ^ (new_n566_ | (~new_n564_ & (new_n569_ | (~new_n571_ & (new_n530_ | new_n570_))))));
  assign new_n865_ = ((~new_n348_ & new_n537_) | (~new_n350_ & new_n533_)) ^ (new_n536_ ^ ((~new_n348_ & new_n533_) | (~new_n350_ & new_n535_)));
  assign new_n866_ = (new_n731_ | (~new_n349_ & ~REG3_REG_17__SCAN_IN) | (new_n349_ & REG3_REG_17__SCAN_IN)) & ~new_n867_ & (STATE_REG_SCAN_IN | ~REG3_REG_17__SCAN_IN) & (~new_n598_ | new_n350_);
  assign new_n867_ = new_n593_ & ((~new_n344_ & new_n584_ & ~new_n262_) | (~new_n359_ & new_n584_ & new_n262_));
  assign new_n868_ = (~new_n694_ | (~new_n869_ & new_n870_)) & (new_n873_ | ~new_n875_ | ((~new_n874_ | ~new_n489_) & ~new_n673_ & (new_n874_ | new_n489_)));
  assign new_n869_ = (new_n468_ | new_n613_ | (new_n499_ & ~new_n425_ & new_n484_ & (new_n605_ | new_n472_))) & ~new_n672_ & (~new_n468_ | (~new_n613_ & (~new_n499_ | new_n425_ | ~new_n484_ | (~new_n605_ & ~new_n472_))));
  assign new_n870_ = new_n871_ & ((~new_n468_ & ~new_n638_ & (new_n617_ | ~new_n639_)) | new_n673_ | (new_n468_ & (new_n638_ | (~new_n617_ & new_n639_))));
  assign new_n871_ = new_n872_ & ((~new_n358_ & DATAI_24_ & (DATAI_23_ | ~new_n660_ | ~new_n680_)) | ~new_n526_ | (new_n660_ & new_n680_ & (new_n358_ | ~DATAI_24_) & (new_n358_ | ~DATAI_23_)));
  assign new_n872_ = (new_n399_ | ~new_n667_) & (~new_n382_ | ~new_n600_) & (new_n374_ | ~new_n644_);
  assign new_n873_ = (new_n489_ | (~new_n399_ & ~new_n401_) | ((~new_n399_ | ~new_n401_) & (~new_n648_ | (new_n647_ & (new_n605_ | new_n472_))))) & new_n652_ & (~new_n489_ | ((new_n399_ | new_n401_) & ((new_n399_ & new_n401_) | (new_n648_ & (~new_n647_ | (~new_n605_ & ~new_n472_))))));
  assign new_n874_ = (new_n399_ | ~new_n401_) & ((new_n399_ & ~new_n401_) | ((new_n378_ | ~new_n382_) & (new_n638_ | (~new_n617_ & new_n639_) | (new_n378_ & ~new_n382_))));
  assign new_n875_ = new_n876_ & ((~new_n489_ & new_n612_ & (~new_n611_ | (~new_n605_ & ~new_n472_))) | new_n643_ | (new_n489_ & (~new_n612_ | (new_n611_ & (new_n605_ | new_n472_)))));
  assign new_n876_ = new_n877_ & ((new_n405_ & (new_n401_ | ~new_n681_ | ~new_n660_ | ~new_n680_)) | ~new_n526_ | (~new_n405_ & ~new_n401_ & new_n681_ & new_n660_ & new_n680_));
  assign new_n877_ = (new_n407_ | ~new_n667_) & (new_n399_ | ~new_n644_) & new_n668_ & (~new_n405_ | ~new_n600_);
  assign new_n878_ = ~new_n879_ & (~new_n713_ | ~ADDR_REG_15__SCAN_IN) & (STATE_REG_SCAN_IN | ~REG3_REG_15__SCAN_IN);
  assign new_n879_ = ~new_n714_ & (((new_n716_ | (new_n342_ & REG2_REG_15__SCAN_IN) | (~new_n342_ & ~REG2_REG_15__SCAN_IN)) & ~new_n685_ & ~new_n262_ & (~new_n716_ | (new_n342_ ^ REG2_REG_15__SCAN_IN))) | (new_n262_ & new_n342_) | ((~new_n342_ | (~new_n880_ & REG1_REG_15__SCAN_IN) | (new_n880_ & ~REG1_REG_15__SCAN_IN)) & new_n685_ & (new_n342_ | (~new_n880_ ^ REG1_REG_15__SCAN_IN))));
  assign new_n880_ = (new_n337_ | ~REG1_REG_14__SCAN_IN) & ((new_n337_ & ~REG1_REG_14__SCAN_IN) | (~new_n704_ & (new_n319_ | ~REG1_REG_13__SCAN_IN)));
  assign new_n881_ = new_n270_ & STATE_REG_SCAN_IN;
endmodule


