// Benchmark "b14_C_sat" written by ABC on Thu Oct 20 19:28:06 2022

module b14_C_sat ( 
    DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_,
    DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_,
    DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_,
    DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_,
    DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_,
    STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN,
    REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN,
    REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN,
    REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN,
    REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN,
    REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN,
    REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN,
    REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN,
    IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN,
    IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN,
    IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN,
    IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN,
    IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN,
    IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN,
    IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN,
    IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN,
    IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN,
    IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN,
    IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, D_REG_1__SCAN_IN,
    D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN,
    D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
    D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
    D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
    D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
    D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
    D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
    D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
    D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
    D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
    REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
    REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
    REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
    REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
    REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
    REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
    REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
    REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
    REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
    REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG1_REG_0__SCAN_IN,
    REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN,
    REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN,
    REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN,
    REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN,
    REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN,
    REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN,
    REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN,
    REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN,
    REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN,
    REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN,
    REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
    REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
    REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
    REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
    REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
    REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
    REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
    REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
    REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
    REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
    REG2_REG_30__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN,
    ADDR_REG_11__SCAN_IN, ADDR_REG_1__SCAN_IN, DATAO_REG_7__SCAN_IN,
    DATAO_REG_10__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_21__SCAN_IN,
    DATAO_REG_22__SCAN_IN, DATAO_REG_26__SCAN_IN, B_REG_SCAN_IN,
    REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
    REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
    REG3_REG_22__SCAN_IN,
    sat  );
  input  DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
    DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
    DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
    DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
    DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
    DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN,
    REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN,
    REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN,
    REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN,
    REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN,
    REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN,
    REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN,
    REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN,
    IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN,
    IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN,
    IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN,
    IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN,
    IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN,
    IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN,
    IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN,
    IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN,
    IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN,
    IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN,
    IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, D_REG_1__SCAN_IN,
    D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN,
    D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
    D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
    D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
    D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
    D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
    D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
    D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
    D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
    D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
    REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
    REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
    REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
    REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
    REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
    REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
    REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
    REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
    REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
    REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG1_REG_0__SCAN_IN,
    REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN,
    REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN,
    REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN,
    REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN,
    REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN,
    REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN,
    REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN,
    REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN,
    REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN,
    REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN,
    REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
    REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
    REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
    REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
    REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
    REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
    REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
    REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
    REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
    REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
    REG2_REG_30__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN,
    ADDR_REG_11__SCAN_IN, ADDR_REG_1__SCAN_IN, DATAO_REG_7__SCAN_IN,
    DATAO_REG_10__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_21__SCAN_IN,
    DATAO_REG_22__SCAN_IN, DATAO_REG_26__SCAN_IN, B_REG_SCAN_IN,
    REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
    REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
    REG3_REG_22__SCAN_IN;
  output sat;
  wire new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_;
  assign sat = ((new_n233_ & new_n673_) | ~new_n555_ | (~new_n233_ & ~new_n673_)) & new_n665_ & ~new_n402_ & new_n657_ & new_n501_ & new_n530_;
  assign new_n233_ = ~new_n388_ & (new_n234_ | ~new_n401_ | ~new_n390_);
  assign new_n234_ = new_n381_ & (new_n375_ | (new_n362_ & (new_n235_ | ~new_n363_ | ~new_n387_)));
  assign new_n235_ = ~new_n347_ & new_n355_ & (~new_n334_ | (~new_n361_ & (new_n356_ | new_n360_) & ((~new_n236_ & new_n330_) | (new_n356_ & new_n360_))));
  assign new_n236_ = new_n300_ & ((~new_n319_ & (new_n296_ | (new_n276_ & (new_n324_ | (~new_n237_ & new_n328_))))) | (~new_n329_ & (~new_n319_ | new_n296_ | (new_n276_ & (new_n324_ | (~new_n237_ & new_n328_))))));
  assign new_n237_ = new_n273_ & (~new_n268_ | ((new_n238_ | (~new_n261_ ^ ~new_n269_)) & ((~new_n267_ & ~new_n269_) | (new_n266_ & ~new_n263_ & new_n269_))));
  assign new_n238_ = (~new_n239_ | new_n251_) & (~new_n250_ | new_n256_);
  assign new_n239_ = ~new_n240_ & ((new_n248_ & (IR_REG_31__SCAN_IN ? ((new_n245_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN) | (IR_REG_21__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN))) : ~IR_REG_21__SCAN_IN)) | (~new_n248_ & ~new_n249_) | (~IR_REG_20__SCAN_IN ^ (new_n245_ | ~IR_REG_31__SCAN_IN)));
  assign new_n240_ = ((IR_REG_25__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & (IR_REG_25__SCAN_IN | IR_REG_24__SCAN_IN | ~new_n243_ | ~new_n244_ | ~new_n241_ | ~new_n242_) & (~IR_REG_25__SCAN_IN | (~IR_REG_24__SCAN_IN & new_n243_ & new_n244_ & new_n241_ & new_n242_)))) & (IR_REG_24__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_24__SCAN_IN ^ (new_n243_ & new_n244_ & new_n241_ & new_n242_))) & (~IR_REG_26__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_25__SCAN_IN & ~IR_REG_24__SCAN_IN & new_n243_ & new_n244_ & new_n241_ & new_n242_)));
  assign new_n241_ = ~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN & ~IR_REG_4__SCAN_IN & ~IR_REG_5__SCAN_IN & ~IR_REG_3__SCAN_IN & ~IR_REG_6__SCAN_IN;
  assign new_n242_ = ~IR_REG_13__SCAN_IN & ~IR_REG_11__SCAN_IN & ~IR_REG_12__SCAN_IN & ~IR_REG_9__SCAN_IN & ~IR_REG_10__SCAN_IN & ~IR_REG_7__SCAN_IN & ~IR_REG_8__SCAN_IN;
  assign new_n243_ = ~IR_REG_22__SCAN_IN & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN;
  assign new_n244_ = ~IR_REG_23__SCAN_IN & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN & ~IR_REG_15__SCAN_IN & ~IR_REG_16__SCAN_IN & ~IR_REG_14__SCAN_IN & ~IR_REG_17__SCAN_IN;
  assign new_n245_ = new_n247_ & new_n246_ & new_n241_ & new_n242_;
  assign new_n246_ = ~IR_REG_15__SCAN_IN & ~IR_REG_16__SCAN_IN & ~IR_REG_14__SCAN_IN & ~IR_REG_17__SCAN_IN;
  assign new_n247_ = ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN;
  assign new_n248_ = IR_REG_19__SCAN_IN ^ ((IR_REG_31__SCAN_IN & (~new_n246_ | ~new_n241_ | ~new_n242_)) | (IR_REG_18__SCAN_IN & IR_REG_31__SCAN_IN));
  assign new_n249_ = (~IR_REG_22__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_22__SCAN_IN & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n247_ & new_n246_ & new_n241_ & new_n242_) | (IR_REG_22__SCAN_IN & (IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n247_ | ~new_n246_ | ~new_n241_ | ~new_n242_)));
  assign new_n250_ = ~new_n240_ & (~IR_REG_31__SCAN_IN | ((~new_n245_ | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN) & (~IR_REG_21__SCAN_IN | (new_n245_ & ~IR_REG_20__SCAN_IN)))) & (IR_REG_21__SCAN_IN | IR_REG_31__SCAN_IN) & (IR_REG_20__SCAN_IN ^ (new_n245_ | ~IR_REG_31__SCAN_IN));
  assign new_n251_ = (~REG2_REG_1__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG3_REG_1__SCAN_IN | ~new_n252_ | new_n255_) & (~REG1_REG_1__SCAN_IN | new_n252_ | new_n255_) & (~REG0_REG_1__SCAN_IN | new_n252_ | ~new_n255_);
  assign new_n252_ = IR_REG_31__SCAN_IN ? (~IR_REG_30__SCAN_IN ^ (new_n254_ & new_n253_ & new_n243_ & new_n244_ & new_n241_ & new_n242_)) : IR_REG_30__SCAN_IN;
  assign new_n253_ = ~IR_REG_25__SCAN_IN & ~IR_REG_26__SCAN_IN & ~IR_REG_24__SCAN_IN & ~IR_REG_27__SCAN_IN;
  assign new_n254_ = ~IR_REG_28__SCAN_IN & ~IR_REG_29__SCAN_IN;
  assign new_n255_ = IR_REG_29__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_28__SCAN_IN & new_n253_ & new_n243_ & new_n244_ & new_n241_ & new_n242_));
  assign new_n256_ = (new_n257_ & ~new_n258_) ? ~new_n260_ : ~DATAI_1_;
  assign new_n257_ = (~IR_REG_28__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_28__SCAN_IN & new_n253_ & new_n243_ & new_n244_ & new_n241_ & new_n242_) | (IR_REG_28__SCAN_IN & (~new_n253_ | ~new_n243_ | ~new_n244_ | ~new_n241_ | ~new_n242_)));
  assign new_n258_ = IR_REG_31__SCAN_IN ? ((~new_n243_ | ~new_n244_ | ~new_n241_ | ~new_n242_ | ~new_n259_ | IR_REG_24__SCAN_IN | IR_REG_27__SCAN_IN) & (~IR_REG_27__SCAN_IN | (new_n259_ & ~IR_REG_24__SCAN_IN & new_n243_ & new_n244_ & new_n241_ & new_n242_))) : IR_REG_27__SCAN_IN;
  assign new_n259_ = ~IR_REG_25__SCAN_IN & ~IR_REG_26__SCAN_IN;
  assign new_n260_ = ~IR_REG_1__SCAN_IN ^ (~IR_REG_0__SCAN_IN | ~IR_REG_31__SCAN_IN);
  assign new_n261_ = (~new_n250_ | new_n251_) & (~new_n262_ | new_n256_);
  assign new_n262_ = ~new_n240_ & ((new_n248_ & (IR_REG_31__SCAN_IN ? ((new_n245_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN) | (IR_REG_21__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN))) : ~IR_REG_21__SCAN_IN)) | (~new_n248_ & ~new_n249_) | (~IR_REG_20__SCAN_IN ^ (new_n245_ | ~IR_REG_31__SCAN_IN)) | (new_n249_ & (IR_REG_31__SCAN_IN ? ((new_n245_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN) | (IR_REG_21__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN))) : ~IR_REG_21__SCAN_IN)));
  assign new_n263_ = (~new_n262_ | new_n264_) & (~new_n250_ | new_n265_);
  assign new_n264_ = (new_n257_ & ~new_n258_) ? ~IR_REG_0__SCAN_IN : ~DATAI_0_;
  assign new_n265_ = (~REG2_REG_0__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG3_REG_0__SCAN_IN | ~new_n252_ | new_n255_) & (~REG1_REG_0__SCAN_IN | new_n252_ | new_n255_) & (~REG0_REG_0__SCAN_IN | new_n252_ | ~new_n255_);
  assign new_n266_ = (~new_n250_ | new_n264_) & (~new_n239_ | new_n265_);
  assign new_n267_ = ((new_n250_ & ~new_n265_) | (new_n262_ & ~new_n264_) | (new_n240_ & REG1_REG_0__SCAN_IN)) & ((new_n240_ & IR_REG_0__SCAN_IN) | (new_n250_ & ~new_n264_) | (new_n239_ & ~new_n265_));
  assign new_n268_ = ((new_n239_ & ~new_n270_) | (new_n250_ & ~new_n271_) | (~new_n269_ & ((new_n250_ & ~new_n270_) | (new_n262_ & ~new_n271_))) | (new_n269_ & (~new_n250_ | new_n270_) & (~new_n262_ | new_n271_))) & ((new_n239_ & ~new_n251_) | (new_n250_ & ~new_n256_) | (~new_n269_ & ((new_n250_ & ~new_n251_) | (new_n262_ & ~new_n256_))) | (new_n269_ & (~new_n250_ | new_n251_) & (~new_n262_ | new_n256_)));
  assign new_n269_ = ((IR_REG_31__SCAN_IN ? ((~new_n245_ | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN) & (~IR_REG_21__SCAN_IN | (new_n245_ & ~IR_REG_20__SCAN_IN))) : IR_REG_21__SCAN_IN) | new_n248_ | new_n249_) & ~new_n240_ & ((~IR_REG_21__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & ((new_n245_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN) | (IR_REG_21__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN)))) | (~IR_REG_20__SCAN_IN ^ (new_n245_ | ~IR_REG_31__SCAN_IN)));
  assign new_n270_ = (~REG2_REG_2__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG3_REG_2__SCAN_IN | ~new_n252_ | new_n255_) & (~REG1_REG_2__SCAN_IN | new_n252_ | new_n255_) & (~REG0_REG_2__SCAN_IN | new_n252_ | ~new_n255_);
  assign new_n271_ = (new_n257_ & ~new_n258_) ? new_n272_ : ~DATAI_2_;
  assign new_n272_ = (~IR_REG_2__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN) | (IR_REG_2__SCAN_IN & (IR_REG_0__SCAN_IN | IR_REG_1__SCAN_IN)));
  assign new_n273_ = (((~new_n239_ | new_n270_) & (~new_n250_ | new_n271_)) | (~new_n269_ ^ ((new_n250_ & ~new_n270_) | (new_n262_ & ~new_n271_)))) & (((~new_n239_ | new_n274_) & (~new_n250_ | new_n275_)) | (~new_n269_ ^ ((new_n250_ & ~new_n274_) | (new_n262_ & ~new_n275_))));
  assign new_n274_ = (~REG1_REG_3__SCAN_IN | new_n252_ | new_n255_) & (~REG0_REG_3__SCAN_IN | new_n252_ | ~new_n255_) & (~REG2_REG_3__SCAN_IN | ~new_n252_ | ~new_n255_) & (REG3_REG_3__SCAN_IN | ~new_n252_ | new_n255_);
  assign new_n275_ = (new_n257_ & ~new_n258_) ? (IR_REG_3__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN))) : ~DATAI_3_;
  assign new_n276_ = ~new_n286_ & ~new_n290_ & ~new_n277_ & ~new_n282_;
  assign new_n277_ = (new_n269_ | ((~new_n250_ | new_n278_) & (~new_n262_ | ~new_n280_))) & (~new_n269_ | (new_n250_ & ~new_n278_) | (new_n262_ & new_n280_)) & (~new_n239_ | new_n278_) & (~new_n250_ | ~new_n280_);
  assign new_n278_ = (~new_n252_ | new_n255_ | (new_n279_ & REG3_REG_7__SCAN_IN & REG3_REG_6__SCAN_IN) | (~REG3_REG_7__SCAN_IN & (~new_n279_ | ~REG3_REG_6__SCAN_IN))) & (~REG1_REG_7__SCAN_IN | new_n252_ | new_n255_) & (~REG2_REG_7__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG0_REG_7__SCAN_IN | new_n252_ | ~new_n255_);
  assign new_n279_ = REG3_REG_5__SCAN_IN & REG3_REG_3__SCAN_IN & REG3_REG_4__SCAN_IN;
  assign new_n280_ = (new_n257_ & ~new_n258_) ? new_n281_ : DATAI_7_;
  assign new_n281_ = IR_REG_31__SCAN_IN ? (~new_n241_ ^ IR_REG_7__SCAN_IN) : IR_REG_7__SCAN_IN;
  assign new_n282_ = (~new_n239_ | new_n283_) & (~new_n250_ | new_n284_) & (new_n269_ | ((~new_n250_ | new_n283_) & (~new_n262_ | new_n284_))) & (~new_n269_ | (new_n250_ & ~new_n283_) | (new_n262_ & ~new_n284_));
  assign new_n283_ = (~REG2_REG_6__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG1_REG_6__SCAN_IN | new_n252_ | new_n255_) & (~REG0_REG_6__SCAN_IN | new_n252_ | ~new_n255_) & (~new_n252_ | new_n255_ | (new_n279_ & REG3_REG_6__SCAN_IN) | (~new_n279_ & ~REG3_REG_6__SCAN_IN));
  assign new_n284_ = (new_n257_ & ~new_n258_) ? new_n285_ : ~DATAI_6_;
  assign new_n285_ = (~IR_REG_6__SCAN_IN | IR_REG_31__SCAN_IN) & ((IR_REG_6__SCAN_IN & (IR_REG_4__SCAN_IN | IR_REG_5__SCAN_IN | IR_REG_3__SCAN_IN | IR_REG_2__SCAN_IN | IR_REG_0__SCAN_IN | IR_REG_1__SCAN_IN)) | ~IR_REG_31__SCAN_IN | (~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN & ~IR_REG_4__SCAN_IN & ~IR_REG_5__SCAN_IN & ~IR_REG_3__SCAN_IN & ~IR_REG_6__SCAN_IN));
  assign new_n286_ = (~new_n239_ | new_n287_) & (~new_n250_ | new_n288_) & (new_n269_ | ((~new_n250_ | new_n287_) & (~new_n262_ | new_n288_))) & (~new_n269_ | (new_n250_ & ~new_n287_) | (new_n262_ & ~new_n288_));
  assign new_n287_ = (~REG2_REG_5__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG1_REG_5__SCAN_IN | new_n252_ | new_n255_) & (~REG0_REG_5__SCAN_IN | new_n252_ | ~new_n255_) & (~new_n252_ | new_n255_ | (REG3_REG_5__SCAN_IN & REG3_REG_3__SCAN_IN & REG3_REG_4__SCAN_IN) | (~REG3_REG_5__SCAN_IN & (~REG3_REG_3__SCAN_IN | ~REG3_REG_4__SCAN_IN)));
  assign new_n288_ = (new_n257_ & ~new_n258_) ? ~new_n289_ : ~DATAI_5_;
  assign new_n289_ = IR_REG_5__SCAN_IN ^ ((IR_REG_31__SCAN_IN & (IR_REG_3__SCAN_IN | IR_REG_2__SCAN_IN | IR_REG_0__SCAN_IN | IR_REG_1__SCAN_IN)) | (IR_REG_4__SCAN_IN & IR_REG_31__SCAN_IN));
  assign new_n290_ = (~new_n239_ | new_n291_) & (~new_n250_ | new_n293_) & (new_n269_ | ((~new_n250_ | new_n291_) & (~new_n262_ | new_n293_))) & (~new_n269_ | (new_n250_ & ~new_n291_) | (new_n262_ & ~new_n293_));
  assign new_n291_ = (~REG2_REG_8__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG1_REG_8__SCAN_IN | new_n252_ | new_n255_) & (~new_n292_ | ~new_n252_ | new_n255_) & (~REG0_REG_8__SCAN_IN | new_n252_ | ~new_n255_);
  assign new_n292_ = REG3_REG_8__SCAN_IN ^ (new_n279_ & REG3_REG_7__SCAN_IN & REG3_REG_6__SCAN_IN);
  assign new_n293_ = (new_n257_ & ~new_n258_) ? new_n294_ : ~DATAI_8_;
  assign new_n294_ = (~IR_REG_8__SCAN_IN | IR_REG_31__SCAN_IN) & ((~new_n295_ & IR_REG_8__SCAN_IN) | ~IR_REG_31__SCAN_IN | (new_n295_ & ~IR_REG_8__SCAN_IN));
  assign new_n295_ = ~IR_REG_7__SCAN_IN & ~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN & ~IR_REG_4__SCAN_IN & ~IR_REG_5__SCAN_IN & ~IR_REG_3__SCAN_IN & ~IR_REG_6__SCAN_IN;
  assign new_n296_ = ~new_n290_ & ((new_n297_ & ~new_n277_ & ~new_n282_) | ~new_n299_ | (~new_n277_ & new_n298_));
  assign new_n297_ = ((new_n239_ & ~new_n287_) | (new_n250_ & ~new_n288_)) & (new_n269_ ^ ((new_n250_ & ~new_n287_) | (new_n262_ & ~new_n288_)));
  assign new_n298_ = ((new_n239_ & ~new_n283_) | (new_n250_ & ~new_n284_)) & (new_n269_ ^ ((new_n250_ & ~new_n283_) | (new_n262_ & ~new_n284_)));
  assign new_n299_ = (((~new_n239_ | new_n291_) & (~new_n250_ | new_n293_)) | (~new_n269_ ^ ((new_n250_ & ~new_n291_) | (new_n262_ & ~new_n293_)))) & ((~new_n269_ ^ ((new_n250_ & ~new_n278_) | (new_n262_ & new_n280_))) | ((~new_n239_ | new_n278_) & (~new_n250_ | ~new_n280_)));
  assign new_n300_ = ~new_n301_ & new_n310_;
  assign new_n301_ = (((~new_n239_ | new_n306_) & (~new_n250_ | new_n308_) & (new_n269_ | ((~new_n250_ | new_n306_) & (~new_n262_ | new_n308_))) & (~new_n269_ | (new_n250_ & ~new_n306_) | (new_n262_ & ~new_n308_))) | (~new_n269_ ^ ((new_n250_ & ~new_n302_) | (new_n262_ & ~new_n304_)))) & (((~new_n239_ | new_n306_) & (~new_n250_ | new_n308_) & (new_n269_ | ((~new_n250_ | new_n306_) & (~new_n262_ | new_n308_))) & (~new_n269_ | (new_n250_ & ~new_n306_) | (new_n262_ & ~new_n308_))) | ((~new_n239_ | new_n302_) & (~new_n250_ | new_n304_)));
  assign new_n302_ = (~REG2_REG_10__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG1_REG_10__SCAN_IN | new_n252_ | new_n255_) & (~new_n303_ | ~new_n252_ | new_n255_) & (~REG0_REG_10__SCAN_IN | new_n252_ | ~new_n255_);
  assign new_n303_ = REG3_REG_10__SCAN_IN ^ (REG3_REG_9__SCAN_IN & REG3_REG_8__SCAN_IN & new_n279_ & REG3_REG_7__SCAN_IN & REG3_REG_6__SCAN_IN);
  assign new_n304_ = (new_n257_ & ~new_n258_) ? new_n305_ : ~DATAI_10_;
  assign new_n305_ = (~IR_REG_10__SCAN_IN | IR_REG_31__SCAN_IN) & ((IR_REG_10__SCAN_IN & (IR_REG_9__SCAN_IN | ~new_n295_ | IR_REG_8__SCAN_IN)) | ~IR_REG_31__SCAN_IN | (~IR_REG_10__SCAN_IN & ~IR_REG_9__SCAN_IN & new_n295_ & ~IR_REG_8__SCAN_IN));
  assign new_n306_ = (~REG2_REG_11__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG1_REG_11__SCAN_IN | new_n252_ | new_n255_) & (~REG0_REG_11__SCAN_IN | new_n252_ | ~new_n255_) & (~new_n252_ | new_n255_ | (new_n307_ & REG3_REG_11__SCAN_IN) | (~new_n307_ & ~REG3_REG_11__SCAN_IN));
  assign new_n307_ = REG3_REG_10__SCAN_IN & REG3_REG_9__SCAN_IN & REG3_REG_8__SCAN_IN & REG3_REG_5__SCAN_IN & REG3_REG_3__SCAN_IN & REG3_REG_4__SCAN_IN & REG3_REG_7__SCAN_IN & REG3_REG_6__SCAN_IN;
  assign new_n308_ = (new_n257_ & ~new_n258_) ? ~new_n309_ : ~DATAI_11_;
  assign new_n309_ = IR_REG_31__SCAN_IN ? (IR_REG_11__SCAN_IN ^ (IR_REG_10__SCAN_IN | IR_REG_9__SCAN_IN | ~new_n295_ | IR_REG_8__SCAN_IN)) : IR_REG_11__SCAN_IN;
  assign new_n310_ = ((new_n239_ & ~new_n314_) | (new_n250_ & ~new_n316_) | (~new_n269_ & ((new_n250_ & ~new_n314_) | (new_n262_ & ~new_n316_))) | (new_n269_ & (~new_n250_ | new_n314_) & (~new_n262_ | new_n316_))) & ((new_n239_ & ~new_n311_) | (new_n250_ & ~new_n312_) | (~new_n269_ & ((new_n250_ & ~new_n311_) | (new_n262_ & ~new_n312_))) | (new_n269_ & (~new_n250_ | new_n311_) & (~new_n262_ | new_n312_)));
  assign new_n311_ = (~REG2_REG_12__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG0_REG_12__SCAN_IN | new_n252_ | ~new_n255_) & (~REG1_REG_12__SCAN_IN | new_n252_ | new_n255_) & (~new_n252_ | new_n255_ | (~REG3_REG_12__SCAN_IN & (~new_n307_ | ~REG3_REG_11__SCAN_IN)) | (REG3_REG_12__SCAN_IN & new_n307_ & REG3_REG_11__SCAN_IN));
  assign new_n312_ = (new_n257_ & ~new_n258_) ? ~new_n313_ : ~DATAI_12_;
  assign new_n313_ = ~IR_REG_12__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_11__SCAN_IN & ~IR_REG_10__SCAN_IN & ~IR_REG_9__SCAN_IN & new_n295_ & ~IR_REG_8__SCAN_IN));
  assign new_n314_ = (~REG2_REG_13__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG1_REG_13__SCAN_IN | new_n252_ | new_n255_) & (~new_n315_ | ~new_n252_ | new_n255_) & (~REG0_REG_13__SCAN_IN | new_n252_ | ~new_n255_);
  assign new_n315_ = REG3_REG_13__SCAN_IN ^ (REG3_REG_12__SCAN_IN & new_n307_ & REG3_REG_11__SCAN_IN);
  assign new_n316_ = (new_n257_ & ~new_n258_) ? ((~IR_REG_13__SCAN_IN | IR_REG_31__SCAN_IN) & (new_n317_ | ~IR_REG_31__SCAN_IN | (IR_REG_13__SCAN_IN & (~new_n318_ | IR_REG_12__SCAN_IN)))) : ~DATAI_13_;
  assign new_n317_ = new_n241_ & new_n242_;
  assign new_n318_ = ~IR_REG_11__SCAN_IN & ~IR_REG_10__SCAN_IN & ~IR_REG_9__SCAN_IN & new_n295_ & ~IR_REG_8__SCAN_IN;
  assign new_n319_ = (~new_n239_ | new_n320_) & (~new_n250_ | new_n322_);
  assign new_n320_ = (~REG2_REG_9__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG0_REG_9__SCAN_IN | new_n252_ | ~new_n255_) & (~new_n321_ | ~new_n252_ | new_n255_) & (~REG1_REG_9__SCAN_IN | new_n252_ | new_n255_);
  assign new_n321_ = REG3_REG_9__SCAN_IN ^ (REG3_REG_8__SCAN_IN & new_n279_ & REG3_REG_7__SCAN_IN & REG3_REG_6__SCAN_IN);
  assign new_n322_ = (new_n257_ & ~new_n258_) ? new_n323_ : ~DATAI_9_;
  assign new_n323_ = IR_REG_9__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (new_n295_ & ~IR_REG_8__SCAN_IN));
  assign new_n324_ = ((new_n239_ & ~new_n325_) | (new_n250_ & ~new_n326_)) & (new_n269_ ^ ((new_n250_ & ~new_n325_) | (new_n262_ & ~new_n326_)));
  assign new_n325_ = (~REG1_REG_4__SCAN_IN | new_n252_ | new_n255_) & (~REG2_REG_4__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG0_REG_4__SCAN_IN | new_n252_ | ~new_n255_) & (~new_n252_ | new_n255_ | (REG3_REG_3__SCAN_IN & REG3_REG_4__SCAN_IN) | (~REG3_REG_3__SCAN_IN & ~REG3_REG_4__SCAN_IN));
  assign new_n326_ = (new_n257_ & ~new_n258_) ? new_n327_ : ~DATAI_4_;
  assign new_n327_ = IR_REG_4__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_3__SCAN_IN & ~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN));
  assign new_n328_ = ((new_n239_ & ~new_n274_) | (new_n250_ & ~new_n275_) | (~new_n269_ & ((new_n250_ & ~new_n274_) | (new_n262_ & ~new_n275_))) | (new_n269_ & (~new_n250_ | new_n274_) & (~new_n262_ | new_n275_))) & ((new_n239_ & ~new_n325_) | (new_n250_ & ~new_n326_) | (~new_n269_ & ((new_n250_ & ~new_n325_) | (new_n262_ & ~new_n326_))) | (new_n269_ & (~new_n250_ | new_n325_) & (~new_n262_ | new_n326_)));
  assign new_n329_ = ~new_n269_ ^ ((new_n250_ & ~new_n320_) | (new_n262_ & ~new_n322_));
  assign new_n330_ = (new_n331_ | ~new_n310_) & ((~new_n269_ ^ ((new_n262_ & ~new_n316_) | (new_n250_ & ~new_n314_))) | ((~new_n250_ | new_n316_) & (~new_n239_ | new_n314_)));
  assign new_n331_ = ~new_n332_ & ~new_n333_ & ((~new_n269_ ^ ((new_n262_ & ~new_n312_) | (new_n250_ & ~new_n311_))) | ((~new_n250_ | new_n312_) & (~new_n239_ | new_n311_)));
  assign new_n332_ = (new_n269_ ^ ((new_n250_ & ~new_n302_) | (new_n262_ & ~new_n304_))) & ((new_n239_ & ~new_n306_) | (new_n250_ & ~new_n308_) | (~new_n269_ & ((new_n250_ & ~new_n306_) | (new_n262_ & ~new_n308_))) | (new_n269_ & (~new_n250_ | new_n306_) & (~new_n262_ | new_n308_))) & ((new_n239_ & ~new_n302_) | (new_n250_ & ~new_n304_));
  assign new_n333_ = ((new_n239_ & ~new_n306_) | (new_n250_ & ~new_n308_)) & (new_n269_ ^ ((new_n250_ & ~new_n306_) | (new_n262_ & ~new_n308_)));
  assign new_n334_ = new_n335_ & ((~new_n269_ & ((new_n250_ & ~new_n345_) | (new_n262_ & ~new_n346_))) | (new_n269_ & (~new_n250_ | new_n345_) & (~new_n262_ | new_n346_)) | (new_n239_ & ~new_n345_) | (new_n250_ & ~new_n346_));
  assign new_n335_ = ((~new_n269_ & ((new_n250_ & ~new_n340_) | (new_n262_ & ~new_n342_))) | (new_n269_ & (~new_n250_ | new_n340_) & (~new_n262_ | new_n342_)) | (new_n239_ & ~new_n340_) | (new_n250_ & ~new_n342_)) & ((~new_n336_ & new_n239_) | (new_n250_ & ~new_n343_) | (~new_n269_ & ((~new_n336_ & new_n250_) | (new_n262_ & ~new_n343_))) | (new_n269_ & (new_n336_ | ~new_n250_) & (~new_n262_ | new_n343_)));
  assign new_n336_ = ~new_n337_ & new_n339_;
  assign new_n337_ = (REG3_REG_17__SCAN_IN | (new_n338_ & REG3_REG_16__SCAN_IN)) & (~REG3_REG_17__SCAN_IN | ~new_n338_ | ~REG3_REG_16__SCAN_IN) & new_n252_ & ~new_n255_;
  assign new_n338_ = REG3_REG_15__SCAN_IN & REG3_REG_14__SCAN_IN & REG3_REG_13__SCAN_IN & REG3_REG_12__SCAN_IN & new_n307_ & REG3_REG_11__SCAN_IN;
  assign new_n339_ = (~REG0_REG_17__SCAN_IN | new_n252_ | ~new_n255_) & (~REG2_REG_17__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG1_REG_17__SCAN_IN | new_n252_ | new_n255_);
  assign new_n340_ = (~REG2_REG_15__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG0_REG_15__SCAN_IN | new_n252_ | ~new_n255_) & (~new_n341_ | ~new_n252_ | new_n255_) & (~REG1_REG_15__SCAN_IN | new_n252_ | new_n255_);
  assign new_n341_ = REG3_REG_15__SCAN_IN ^ (REG3_REG_14__SCAN_IN & REG3_REG_13__SCAN_IN & REG3_REG_12__SCAN_IN & new_n307_ & REG3_REG_11__SCAN_IN);
  assign new_n342_ = (new_n257_ & ~new_n258_) ? ((~IR_REG_15__SCAN_IN & (~IR_REG_31__SCAN_IN | (new_n317_ & ~IR_REG_14__SCAN_IN))) | (IR_REG_15__SCAN_IN & IR_REG_31__SCAN_IN & (~new_n317_ | IR_REG_14__SCAN_IN))) : ~DATAI_15_;
  assign new_n343_ = (new_n257_ & ~new_n258_) ? ~new_n344_ : ~DATAI_17_;
  assign new_n344_ = ~IR_REG_17__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_15__SCAN_IN & ~IR_REG_16__SCAN_IN & ~IR_REG_14__SCAN_IN & new_n241_ & new_n242_));
  assign new_n345_ = ((~new_n338_ & ~REG3_REG_16__SCAN_IN) | (new_n338_ & REG3_REG_16__SCAN_IN) | ~new_n252_ | new_n255_) & (~REG0_REG_16__SCAN_IN | new_n252_ | ~new_n255_) & (~REG1_REG_16__SCAN_IN | new_n252_ | new_n255_) & (~REG2_REG_16__SCAN_IN | ~new_n252_ | ~new_n255_);
  assign new_n346_ = (new_n257_ & ~new_n258_) ? (~IR_REG_16__SCAN_IN ^ ((IR_REG_15__SCAN_IN & IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & (~new_n317_ | IR_REG_14__SCAN_IN)))) : ~DATAI_16_;
  assign new_n347_ = ~new_n348_ & ~new_n354_;
  assign new_n348_ = (~new_n239_ | new_n352_) & (new_n349_ | ~new_n250_);
  assign new_n349_ = new_n351_ ? (IR_REG_18__SCAN_IN ^ (new_n350_ | ~IR_REG_31__SCAN_IN)) : ~DATAI_18_;
  assign new_n350_ = new_n317_ & new_n246_;
  assign new_n351_ = new_n257_ & ~new_n258_;
  assign new_n352_ = (~new_n252_ | new_n255_ | (new_n353_ & REG3_REG_18__SCAN_IN) | (~new_n353_ & ~REG3_REG_18__SCAN_IN)) & (~REG1_REG_18__SCAN_IN | new_n252_ | new_n255_) & (~REG2_REG_18__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG0_REG_18__SCAN_IN | new_n252_ | ~new_n255_);
  assign new_n353_ = REG3_REG_17__SCAN_IN & REG3_REG_16__SCAN_IN & REG3_REG_15__SCAN_IN & REG3_REG_14__SCAN_IN & REG3_REG_13__SCAN_IN & REG3_REG_12__SCAN_IN & new_n307_ & REG3_REG_11__SCAN_IN;
  assign new_n354_ = ~new_n269_ ^ ((new_n250_ & ~new_n352_) | (~new_n349_ & new_n262_));
  assign new_n355_ = (((new_n336_ | ~new_n239_) & (~new_n250_ | new_n343_)) | (~new_n269_ ^ ((~new_n336_ & new_n250_) | (new_n262_ & ~new_n343_)))) & (((new_n336_ | ~new_n239_) & (~new_n250_ | new_n343_) & (new_n269_ | ((new_n336_ | ~new_n250_) & (~new_n262_ | new_n343_))) & (~new_n269_ | (~new_n336_ & new_n250_) | (new_n262_ & ~new_n343_))) | (~new_n269_ ^ ((new_n250_ & ~new_n345_) | (new_n262_ & ~new_n346_))) | ((~new_n239_ | new_n345_) & (~new_n250_ | new_n346_)));
  assign new_n356_ = (new_n357_ | ~new_n239_) & (new_n359_ | ~new_n250_);
  assign new_n357_ = (~REG2_REG_14__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG1_REG_14__SCAN_IN | new_n252_ | new_n255_) & (~new_n358_ | ~new_n252_ | new_n255_) & (~REG0_REG_14__SCAN_IN | new_n252_ | ~new_n255_);
  assign new_n358_ = REG3_REG_14__SCAN_IN ^ (REG3_REG_13__SCAN_IN & REG3_REG_12__SCAN_IN & new_n307_ & REG3_REG_11__SCAN_IN);
  assign new_n359_ = (new_n257_ & ~new_n258_) ? (IR_REG_14__SCAN_IN ^ (new_n317_ | ~IR_REG_31__SCAN_IN)) : ~DATAI_14_;
  assign new_n360_ = ~new_n269_ ^ ((~new_n359_ & new_n262_) | (~new_n357_ & new_n250_));
  assign new_n361_ = ((new_n239_ & ~new_n340_) | (new_n250_ & ~new_n342_)) & (new_n269_ ^ ((new_n250_ & ~new_n340_) | (new_n262_ & ~new_n342_)));
  assign new_n362_ = (~new_n363_ | new_n372_) & ((~new_n269_ ^ ((new_n262_ & new_n371_) | (~new_n364_ & new_n250_))) | ((new_n364_ | ~new_n239_) & (~new_n250_ | ~new_n371_)));
  assign new_n363_ = ((~new_n269_ & ((~new_n364_ & new_n250_) | (new_n262_ & new_n371_))) | (new_n269_ & (new_n364_ | ~new_n250_) & (~new_n262_ | ~new_n371_)) | (~new_n364_ & new_n239_) | (new_n250_ & new_n371_)) & ((new_n370_ & new_n250_) | (~new_n368_ & new_n239_) | (~new_n269_ & ((~new_n368_ & new_n250_) | (new_n370_ & new_n262_))) | (new_n269_ & (new_n368_ | ~new_n250_) & (~new_n370_ | ~new_n262_)));
  assign new_n364_ = new_n367_ & (~new_n365_ | ~new_n366_);
  assign new_n365_ = new_n252_ & ~new_n255_;
  assign new_n366_ = REG3_REG_21__SCAN_IN ^ (REG3_REG_20__SCAN_IN & REG3_REG_19__SCAN_IN & new_n353_ & REG3_REG_18__SCAN_IN);
  assign new_n367_ = (~REG0_REG_21__SCAN_IN | new_n252_ | ~new_n255_) & (~REG2_REG_21__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG1_REG_21__SCAN_IN | new_n252_ | new_n255_);
  assign new_n368_ = (~new_n369_ | ~new_n252_ | new_n255_) & (~REG0_REG_20__SCAN_IN | new_n252_ | ~new_n255_) & (~REG1_REG_20__SCAN_IN | new_n252_ | new_n255_) & (~REG2_REG_20__SCAN_IN | ~new_n252_ | ~new_n255_);
  assign new_n369_ = REG3_REG_20__SCAN_IN ^ (REG3_REG_19__SCAN_IN & new_n353_ & REG3_REG_18__SCAN_IN);
  assign new_n370_ = ~new_n351_ & DATAI_20_;
  assign new_n371_ = DATAI_21_ & (~new_n257_ | new_n258_);
  assign new_n372_ = (((~new_n370_ | ~new_n250_) & (new_n368_ | ~new_n239_)) | (~new_n269_ ^ ((~new_n368_ & new_n250_) | (new_n370_ & new_n262_)))) & (((~new_n239_ | new_n374_) & (new_n373_ | ~new_n250_)) | (~new_n269_ ^ ((new_n250_ & ~new_n374_) | (~new_n373_ & new_n262_))));
  assign new_n373_ = new_n351_ ? ~new_n248_ : ~DATAI_19_;
  assign new_n374_ = ((~REG3_REG_19__SCAN_IN & (~new_n353_ | ~REG3_REG_18__SCAN_IN)) | ~new_n252_ | new_n255_ | (REG3_REG_19__SCAN_IN & new_n353_ & REG3_REG_18__SCAN_IN)) & (~REG1_REG_19__SCAN_IN | new_n252_ | new_n255_) & (~REG2_REG_19__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG0_REG_19__SCAN_IN | new_n252_ | ~new_n255_);
  assign new_n375_ = new_n376_ & (~new_n380_ | ~new_n250_) & (new_n377_ | ~new_n239_);
  assign new_n376_ = ~new_n269_ ^ ((new_n380_ & new_n262_) | (~new_n377_ & new_n250_));
  assign new_n377_ = new_n379_ & (~new_n365_ | ~new_n378_);
  assign new_n378_ = REG3_REG_22__SCAN_IN ^ (REG3_REG_21__SCAN_IN & REG3_REG_20__SCAN_IN & REG3_REG_19__SCAN_IN & new_n353_ & REG3_REG_18__SCAN_IN);
  assign new_n379_ = (~REG1_REG_22__SCAN_IN | new_n252_ | new_n255_) & (~REG2_REG_22__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG0_REG_22__SCAN_IN | new_n252_ | ~new_n255_);
  assign new_n380_ = ~new_n351_ & DATAI_22_;
  assign new_n381_ = (((new_n377_ | ~new_n239_) & (~new_n380_ | ~new_n250_)) | (~new_n269_ ^ ((new_n380_ & new_n262_) | (~new_n377_ & new_n250_)))) & (((~new_n386_ | ~new_n250_) & (new_n382_ | ~new_n239_)) | (~new_n269_ ^ ((new_n386_ & new_n262_) | (~new_n382_ & new_n250_))));
  assign new_n382_ = new_n385_ & (~new_n383_ | ~new_n365_);
  assign new_n383_ = REG3_REG_23__SCAN_IN ^ (REG3_REG_22__SCAN_IN & REG3_REG_21__SCAN_IN & new_n384_ & REG3_REG_20__SCAN_IN);
  assign new_n384_ = REG3_REG_19__SCAN_IN & new_n353_ & REG3_REG_18__SCAN_IN;
  assign new_n385_ = (~REG0_REG_23__SCAN_IN | new_n252_ | ~new_n255_) & (~REG2_REG_23__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG1_REG_23__SCAN_IN | new_n252_ | new_n255_);
  assign new_n386_ = ~new_n351_ & DATAI_23_;
  assign new_n387_ = ((new_n239_ & ~new_n374_) | (~new_n373_ & new_n250_) | (~new_n269_ & ((new_n250_ & ~new_n374_) | (~new_n373_ & new_n262_))) | (new_n269_ & (~new_n250_ | new_n374_) & (new_n373_ | ~new_n262_))) & ((new_n239_ & ~new_n352_) | (~new_n349_ & new_n250_) | (~new_n269_ & ((new_n250_ & ~new_n352_) | (~new_n349_ & new_n262_))) | (new_n269_ & (~new_n250_ | new_n352_) & (new_n349_ | ~new_n262_)));
  assign new_n388_ = ((new_n393_ & new_n250_) | (~new_n391_ & new_n239_) | (~new_n269_ & ((new_n393_ & new_n262_) | (~new_n391_ & new_n250_))) | (new_n269_ & (~new_n393_ | ~new_n262_) & (new_n391_ | ~new_n250_))) & (new_n389_ | new_n400_ | (((new_n393_ & new_n250_) | (~new_n391_ & new_n239_)) & (new_n269_ ^ ((new_n393_ & new_n262_) | (~new_n391_ & new_n250_)))));
  assign new_n389_ = new_n390_ & ((new_n399_ & new_n250_) | (~new_n396_ & new_n239_)) & (new_n269_ ^ ((~new_n396_ & new_n250_) | (new_n399_ & new_n262_)));
  assign new_n390_ = ((new_n395_ & new_n250_) | (~new_n394_ & new_n239_) | (~new_n269_ & ((new_n395_ & new_n262_) | (~new_n394_ & new_n250_))) | (new_n269_ & (~new_n395_ | ~new_n262_) & (new_n394_ | ~new_n250_))) & ((~new_n269_ & ((new_n393_ & new_n262_) | (~new_n391_ & new_n250_))) | (new_n269_ & (~new_n393_ | ~new_n262_) & (new_n391_ | ~new_n250_)) | (new_n393_ & new_n250_) | (~new_n391_ & new_n239_));
  assign new_n391_ = ((REG3_REG_26__SCAN_IN & new_n392_ & REG3_REG_25__SCAN_IN) | ~new_n252_ | new_n255_ | (~REG3_REG_26__SCAN_IN & (~new_n392_ | ~REG3_REG_25__SCAN_IN))) & (~REG1_REG_26__SCAN_IN | new_n252_ | new_n255_) & (~REG2_REG_26__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG0_REG_26__SCAN_IN | new_n252_ | ~new_n255_);
  assign new_n392_ = REG3_REG_24__SCAN_IN & REG3_REG_23__SCAN_IN & REG3_REG_22__SCAN_IN & REG3_REG_21__SCAN_IN & REG3_REG_20__SCAN_IN & REG3_REG_19__SCAN_IN & new_n353_ & REG3_REG_18__SCAN_IN;
  assign new_n393_ = ~new_n351_ & DATAI_26_;
  assign new_n394_ = ((~new_n392_ & ~REG3_REG_25__SCAN_IN) | ~new_n252_ | new_n255_ | (new_n392_ & REG3_REG_25__SCAN_IN)) & (~REG0_REG_25__SCAN_IN | new_n252_ | ~new_n255_) & (~REG1_REG_25__SCAN_IN | new_n252_ | new_n255_) & (~REG2_REG_25__SCAN_IN | ~new_n252_ | ~new_n255_);
  assign new_n395_ = ~new_n351_ & DATAI_25_;
  assign new_n396_ = new_n398_ & ((~REG3_REG_24__SCAN_IN & (~new_n397_ | ~REG3_REG_23__SCAN_IN)) | ~new_n365_ | (REG3_REG_24__SCAN_IN & new_n397_ & REG3_REG_23__SCAN_IN));
  assign new_n397_ = REG3_REG_22__SCAN_IN & REG3_REG_21__SCAN_IN & new_n384_ & REG3_REG_20__SCAN_IN;
  assign new_n398_ = (~REG0_REG_24__SCAN_IN | new_n252_ | ~new_n255_) & (~REG2_REG_24__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG1_REG_24__SCAN_IN | new_n252_ | new_n255_);
  assign new_n399_ = ~new_n351_ & DATAI_24_;
  assign new_n400_ = ((new_n395_ & new_n250_) | (~new_n394_ & new_n239_)) & (new_n269_ ^ ((new_n395_ & new_n262_) | (~new_n394_ & new_n250_)));
  assign new_n401_ = ((~new_n382_ & new_n239_) | (new_n386_ & new_n250_) | (~new_n269_ & ((new_n386_ & new_n262_) | (~new_n382_ & new_n250_))) | (new_n269_ & (~new_n386_ | ~new_n262_) & (new_n382_ | ~new_n250_))) & ((new_n399_ & new_n250_) | (~new_n396_ & new_n239_) | (~new_n269_ & ((new_n399_ & new_n262_) | (~new_n396_ & new_n250_))) | (new_n269_ & (~new_n399_ | ~new_n262_) & (new_n396_ | ~new_n250_)));
  assign new_n402_ = (~new_n474_ | (~new_n403_ & new_n438_)) & ~new_n472_ & new_n494_ & ((new_n489_ & ~new_n435_) | ~new_n500_ | (~new_n489_ & new_n435_));
  assign new_n403_ = ((~new_n433_ & new_n435_) | (new_n433_ & ~new_n435_) | (new_n431_ & ~new_n437_) | (new_n404_ & (new_n431_ | ~new_n437_))) & ~new_n436_ & (((~new_n431_ | new_n437_) & (~new_n404_ | (~new_n431_ & new_n437_))) | (new_n433_ ^ ~new_n435_));
  assign new_n404_ = new_n430_ & (~new_n427_ | (~new_n405_ & ((new_n377_ & ~new_n380_) | (~new_n406_ & new_n424_ & (new_n377_ | ~new_n380_)))));
  assign new_n405_ = ~new_n382_ & new_n386_;
  assign new_n406_ = new_n407_ & new_n420_ & (~new_n418_ | (new_n416_ & (new_n421_ | (new_n423_ & (~new_n409_ | new_n422_)))));
  assign new_n407_ = ~new_n408_ & (~new_n349_ | ~new_n352_) & (~new_n368_ | new_n370_) & (~new_n373_ | ~new_n374_);
  assign new_n408_ = ~new_n371_ & new_n367_ & (~new_n365_ | ~new_n366_);
  assign new_n409_ = (new_n291_ | new_n293_) & ((new_n291_ & new_n293_) | (new_n415_ & (~new_n414_ | (~new_n410_ & ~new_n413_ & (~new_n411_ | ~new_n412_)))));
  assign new_n410_ = ((~new_n274_ & ~new_n275_) | (~new_n270_ & ~new_n271_)) & (~new_n274_ | ~new_n275_) & (~new_n325_ | ~new_n326_) & (~new_n287_ | ~new_n288_);
  assign new_n411_ = (~new_n251_ | ~new_n256_) & ((~new_n264_ & ~new_n265_) | (~new_n251_ & ~new_n256_));
  assign new_n412_ = (~new_n325_ | ~new_n326_) & (~new_n287_ | ~new_n288_) & (~new_n270_ | ~new_n271_) & (~new_n274_ | ~new_n275_);
  assign new_n413_ = (~new_n287_ | ~new_n288_) & ((~new_n287_ & ~new_n288_) | (~new_n325_ & ~new_n326_));
  assign new_n414_ = (~new_n283_ | ~new_n284_) & (~new_n278_ | new_n280_);
  assign new_n415_ = (new_n278_ | ~new_n280_) & (new_n283_ | new_n284_ | (new_n278_ & ~new_n280_));
  assign new_n416_ = new_n417_ & (~new_n311_ | ~new_n312_) & (~new_n314_ | ~new_n316_);
  assign new_n417_ = (~new_n306_ | ~new_n308_) & (~new_n340_ | ~new_n342_) & (~new_n357_ | ~new_n359_);
  assign new_n418_ = (new_n340_ | new_n342_) & (new_n419_ | (new_n357_ & new_n359_) | (new_n340_ & new_n342_));
  assign new_n419_ = (((new_n311_ | new_n312_) & (new_n306_ | new_n308_)) | (new_n311_ & new_n312_) | (new_n314_ & new_n316_)) & (new_n357_ | new_n359_) & (new_n314_ | new_n316_);
  assign new_n420_ = (~new_n336_ | ~new_n343_) & (~new_n345_ | ~new_n346_);
  assign new_n421_ = ~new_n302_ & ~new_n304_;
  assign new_n422_ = ~new_n320_ & ~new_n322_;
  assign new_n423_ = (~new_n302_ | ~new_n304_) & (~new_n320_ | ~new_n322_);
  assign new_n424_ = ~new_n425_ & (~new_n407_ | new_n426_) & (new_n364_ | ~new_n371_);
  assign new_n425_ = ~new_n408_ & ((~new_n368_ & new_n370_) | (~new_n373_ & ~new_n374_ & (~new_n368_ | new_n370_)) | ((~new_n368_ | new_n370_) & (~new_n373_ | ~new_n374_) & ~new_n349_ & ~new_n352_));
  assign new_n426_ = (new_n336_ | new_n343_) & (new_n345_ | new_n346_ | (new_n336_ & new_n343_));
  assign new_n427_ = new_n428_ & ~new_n429_ & (~new_n391_ | new_n393_);
  assign new_n428_ = (new_n399_ | ~new_n398_ | ((REG3_REG_24__SCAN_IN | (new_n397_ & REG3_REG_23__SCAN_IN)) & new_n365_ & (~REG3_REG_24__SCAN_IN | ~new_n397_ | ~REG3_REG_23__SCAN_IN))) & (new_n386_ | ~new_n385_ | (new_n365_ & (~new_n397_ | ~REG3_REG_23__SCAN_IN) & (new_n397_ | REG3_REG_23__SCAN_IN)));
  assign new_n429_ = new_n394_ & ~new_n395_;
  assign new_n430_ = (new_n396_ | ~new_n399_ | (new_n391_ & ~new_n393_) | (new_n394_ & ~new_n395_)) & (new_n391_ | ~new_n393_) & ((new_n391_ & ~new_n393_) | new_n394_ | ~new_n395_);
  assign new_n431_ = (~new_n432_ | ~new_n252_ | new_n255_) & (~REG2_REG_27__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG0_REG_27__SCAN_IN | new_n252_ | ~new_n255_) & (~REG1_REG_27__SCAN_IN | new_n252_ | new_n255_);
  assign new_n432_ = REG3_REG_27__SCAN_IN ^ (REG3_REG_26__SCAN_IN & new_n392_ & REG3_REG_25__SCAN_IN);
  assign new_n433_ = (~REG0_REG_28__SCAN_IN | new_n252_ | ~new_n255_) & (~REG1_REG_28__SCAN_IN | new_n252_ | new_n255_) & (~REG2_REG_28__SCAN_IN | ~new_n252_ | ~new_n255_) & (~new_n252_ | new_n255_ | (~new_n434_ & ~REG3_REG_28__SCAN_IN) | (new_n434_ & REG3_REG_28__SCAN_IN));
  assign new_n434_ = REG3_REG_27__SCAN_IN & REG3_REG_26__SCAN_IN & new_n392_ & REG3_REG_25__SCAN_IN;
  assign new_n435_ = ~new_n351_ & DATAI_28_;
  assign new_n436_ = (((IR_REG_31__SCAN_IN ? ((~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN) | (IR_REG_21__SCAN_IN & (IR_REG_20__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN))) : ~IR_REG_21__SCAN_IN) & (~IR_REG_22__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_22__SCAN_IN & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN) | (IR_REG_22__SCAN_IN & (IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN)))) | ((~IR_REG_31__SCAN_IN | ((IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN) & (~IR_REG_21__SCAN_IN | (~IR_REG_20__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN)))) & (IR_REG_21__SCAN_IN | IR_REG_31__SCAN_IN) & ((IR_REG_22__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & (IR_REG_22__SCAN_IN | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN) & (~IR_REG_22__SCAN_IN | (~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN))))) | (~IR_REG_20__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN))) | (IR_REG_19__SCAN_IN ^ ((~new_n350_ & IR_REG_31__SCAN_IN) | (IR_REG_18__SCAN_IN & IR_REG_31__SCAN_IN)))) & ((~IR_REG_20__SCAN_IN & (~IR_REG_31__SCAN_IN | (new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN))) | (IR_REG_20__SCAN_IN & IR_REG_31__SCAN_IN & (~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN)) | ((~IR_REG_22__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_22__SCAN_IN & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN) | (IR_REG_22__SCAN_IN & (IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN)))) | (IR_REG_19__SCAN_IN ^ ((~new_n350_ & IR_REG_31__SCAN_IN) | (IR_REG_18__SCAN_IN & IR_REG_31__SCAN_IN))));
  assign new_n437_ = DATAI_27_ & (~new_n257_ | new_n258_);
  assign new_n438_ = (new_n431_ | ~new_n468_) & ((~new_n439_ & (~new_n433_ | new_n435_) & (new_n433_ | ~new_n435_)) | new_n470_ | (new_n439_ & (~new_n433_ ^ ~new_n435_)));
  assign new_n439_ = ~new_n440_ & (~new_n465_ | (~new_n466_ & (new_n467_ | (new_n464_ & (~new_n462_ | (new_n441_ & new_n461_))))));
  assign new_n440_ = new_n431_ & new_n437_;
  assign new_n441_ = ~new_n442_ & (~new_n460_ | (new_n459_ & (new_n443_ | ~new_n457_ | (new_n455_ & (new_n444_ | ~new_n453_)))));
  assign new_n442_ = new_n368_ & new_n370_;
  assign new_n443_ = new_n349_ & ~new_n352_;
  assign new_n444_ = new_n451_ & new_n452_ & ((new_n448_ & ~new_n445_ & new_n446_) | ~new_n450_ | (new_n447_ & ~new_n449_));
  assign new_n445_ = ((new_n270_ & ~new_n271_) | ((~new_n256_ | (new_n251_ & ~new_n264_ & new_n265_)) & (new_n251_ | (~new_n264_ & new_n265_)))) & (new_n274_ | ~new_n275_) & (new_n270_ | ~new_n271_);
  assign new_n446_ = (~new_n325_ | new_n326_) & (~new_n274_ | new_n275_);
  assign new_n447_ = (~new_n278_ | ~new_n280_) & (~new_n283_ | new_n284_) & (~new_n291_ | new_n293_);
  assign new_n448_ = (~new_n287_ | new_n288_) & (~new_n278_ | ~new_n280_) & (~new_n291_ | new_n293_) & (~new_n283_ | new_n284_);
  assign new_n449_ = (new_n325_ | ~new_n326_ | (new_n287_ & ~new_n288_)) & (new_n283_ | ~new_n284_) & (new_n287_ | ~new_n288_);
  assign new_n450_ = (new_n291_ | ~new_n293_) & (new_n278_ | new_n280_ | (new_n291_ & ~new_n293_));
  assign new_n451_ = (~new_n302_ | new_n304_) & (~new_n306_ | new_n308_);
  assign new_n452_ = (~new_n320_ | new_n322_) & (~new_n311_ | new_n312_) & (~new_n314_ | new_n316_);
  assign new_n453_ = (new_n314_ | ~new_n316_) & ((new_n314_ & ~new_n316_) | (new_n311_ & ~new_n312_) | (~new_n454_ & (new_n306_ | ~new_n308_) & (new_n311_ | ~new_n312_)));
  assign new_n454_ = ((~new_n320_ & new_n322_) | (~new_n302_ & new_n304_)) & (~new_n302_ | new_n304_) & (~new_n306_ | new_n308_);
  assign new_n455_ = new_n456_ & (~new_n357_ | new_n359_) & (~new_n340_ | new_n342_);
  assign new_n456_ = (~new_n345_ | new_n346_) & (new_n343_ | new_n337_ | ~new_n339_);
  assign new_n457_ = (~new_n456_ | new_n458_) & (new_n336_ | ~new_n343_);
  assign new_n458_ = (new_n340_ | ~new_n342_) & (new_n345_ | ~new_n346_) & ((new_n345_ & ~new_n346_) | new_n357_ | ~new_n359_ | (new_n340_ & ~new_n342_));
  assign new_n459_ = (new_n349_ | ~new_n352_) & (new_n373_ | ~new_n374_);
  assign new_n460_ = (new_n368_ | new_n370_) & (~new_n373_ | new_n374_);
  assign new_n461_ = (~new_n382_ | ~new_n386_) & (~new_n377_ | ~new_n380_) & (~new_n364_ | ~new_n371_);
  assign new_n462_ = new_n463_ & (((new_n377_ | new_n380_) & (new_n364_ | new_n371_)) | (new_n382_ & new_n386_) | (new_n377_ & new_n380_));
  assign new_n463_ = (new_n386_ | (new_n385_ & (~new_n365_ | (new_n397_ & REG3_REG_23__SCAN_IN) | (~new_n397_ & ~REG3_REG_23__SCAN_IN)))) & (new_n399_ | (new_n398_ & ((~REG3_REG_24__SCAN_IN & (~new_n397_ | ~REG3_REG_23__SCAN_IN)) | ~new_n365_ | (REG3_REG_24__SCAN_IN & new_n397_ & REG3_REG_23__SCAN_IN))));
  assign new_n464_ = (~new_n396_ | ~new_n399_) & (~new_n394_ | ~new_n395_);
  assign new_n465_ = (new_n391_ | new_n393_) & (new_n431_ | new_n437_);
  assign new_n466_ = new_n391_ & new_n393_;
  assign new_n467_ = ~new_n394_ & ~new_n395_;
  assign new_n468_ = ~new_n257_ & new_n469_;
  assign new_n469_ = ((IR_REG_22__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & (IR_REG_22__SCAN_IN | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n247_ | ~new_n246_ | ~new_n241_ | ~new_n242_) & (~IR_REG_22__SCAN_IN | (~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n247_ & new_n246_ & new_n241_ & new_n242_)))) & (~IR_REG_31__SCAN_IN | ((IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n247_ | ~new_n246_ | ~new_n241_ | ~new_n242_) & (~IR_REG_21__SCAN_IN | (~IR_REG_20__SCAN_IN & new_n247_ & new_n246_ & new_n241_ & new_n242_)))) & (IR_REG_21__SCAN_IN | IR_REG_31__SCAN_IN);
  assign new_n470_ = (~new_n248_ | new_n249_) & (~new_n471_ | (~IR_REG_21__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & ((new_n245_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN) | (IR_REG_21__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN)))));
  assign new_n471_ = ~IR_REG_20__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (new_n247_ & new_n246_ & new_n241_ & new_n242_));
  assign new_n472_ = ((~new_n433_ & new_n435_) | (new_n433_ & ~new_n435_) | (new_n431_ & ~new_n437_) | (new_n404_ & (new_n431_ | ~new_n437_))) & new_n473_ & (((~new_n431_ | new_n437_) & (~new_n404_ | (~new_n431_ & new_n437_))) | (new_n433_ ^ ~new_n435_));
  assign new_n473_ = new_n474_ & (~IR_REG_19__SCAN_IN | ((new_n350_ | ~IR_REG_31__SCAN_IN) & (~IR_REG_18__SCAN_IN | ~IR_REG_31__SCAN_IN))) & (IR_REG_19__SCAN_IN | (~new_n350_ & IR_REG_31__SCAN_IN) | (IR_REG_18__SCAN_IN & IR_REG_31__SCAN_IN)) & (IR_REG_21__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | ((IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN) & (~IR_REG_21__SCAN_IN | (~IR_REG_20__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN)))) & (IR_REG_20__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN)));
  assign new_n474_ = new_n485_ & (new_n487_ | (new_n479_ & ~new_n475_ & ~new_n488_));
  assign new_n475_ = (new_n477_ | ~new_n478_) & (D_REG_0__SCAN_IN | (new_n476_ & ~new_n477_ & B_REG_SCAN_IN) | new_n478_ | (new_n477_ & ~B_REG_SCAN_IN));
  assign new_n476_ = (~IR_REG_25__SCAN_IN | IR_REG_31__SCAN_IN) & ((IR_REG_25__SCAN_IN & (IR_REG_24__SCAN_IN | ~new_n243_ | ~new_n244_ | ~new_n241_ | ~new_n242_)) | ~IR_REG_31__SCAN_IN | (~IR_REG_25__SCAN_IN & ~IR_REG_24__SCAN_IN & new_n243_ & new_n244_ & new_n241_ & new_n242_));
  assign new_n477_ = IR_REG_31__SCAN_IN ? (~IR_REG_24__SCAN_IN ^ (new_n243_ & new_n244_ & new_n241_ & new_n242_)) : IR_REG_24__SCAN_IN;
  assign new_n478_ = IR_REG_26__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_25__SCAN_IN & ~IR_REG_24__SCAN_IN & new_n243_ & new_n244_ & new_n241_ & new_n242_));
  assign new_n479_ = (new_n480_ | (new_n476_ & ~new_n477_ & B_REG_SCAN_IN) | new_n478_ | (new_n477_ & ~B_REG_SCAN_IN)) & (~new_n476_ | ~new_n478_) & (D_REG_1__SCAN_IN | (new_n476_ & ~new_n477_ & B_REG_SCAN_IN) | new_n478_ | (new_n477_ & ~B_REG_SCAN_IN));
  assign new_n480_ = new_n483_ & new_n484_ & new_n481_ & new_n482_;
  assign new_n481_ = ~D_REG_18__SCAN_IN & ~D_REG_19__SCAN_IN & ~D_REG_16__SCAN_IN & ~D_REG_17__SCAN_IN & ~D_REG_20__SCAN_IN & ~D_REG_21__SCAN_IN & ~D_REG_22__SCAN_IN & ~D_REG_23__SCAN_IN;
  assign new_n482_ = ~D_REG_26__SCAN_IN & ~D_REG_27__SCAN_IN & ~D_REG_24__SCAN_IN & ~D_REG_25__SCAN_IN & ~D_REG_28__SCAN_IN & ~D_REG_29__SCAN_IN & ~D_REG_30__SCAN_IN & ~D_REG_31__SCAN_IN;
  assign new_n483_ = ~D_REG_4__SCAN_IN & ~D_REG_8__SCAN_IN & ~D_REG_2__SCAN_IN & ~D_REG_3__SCAN_IN & ~D_REG_5__SCAN_IN & ~D_REG_6__SCAN_IN;
  assign new_n484_ = ~D_REG_10__SCAN_IN & ~D_REG_11__SCAN_IN & ~D_REG_7__SCAN_IN & ~D_REG_9__SCAN_IN & ~D_REG_12__SCAN_IN & ~D_REG_13__SCAN_IN & ~D_REG_14__SCAN_IN & ~D_REG_15__SCAN_IN;
  assign new_n485_ = STATE_REG_SCAN_IN & ~new_n240_ & ~new_n486_;
  assign new_n486_ = (~IR_REG_23__SCAN_IN | ~IR_REG_31__SCAN_IN | (new_n243_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN & new_n246_ & new_n241_ & new_n242_)) & (IR_REG_23__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | ~new_n241_ | ~new_n242_ | ~new_n243_ | ~new_n246_ | IR_REG_23__SCAN_IN | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN);
  assign new_n487_ = (~IR_REG_22__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (new_n245_ & ~IR_REG_22__SCAN_IN & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN) | (IR_REG_22__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN))) & (IR_REG_20__SCAN_IN ^ (new_n245_ | ~IR_REG_31__SCAN_IN)) & new_n248_ & (IR_REG_31__SCAN_IN ? ((new_n245_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN) | (IR_REG_21__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN))) : ~IR_REG_21__SCAN_IN);
  assign new_n488_ = new_n469_ & (new_n248_ | new_n471_);
  assign new_n489_ = ~new_n437_ & ~new_n393_ & ~new_n395_ & ~new_n399_ & new_n490_ & ~new_n386_;
  assign new_n490_ = ~new_n380_ & ~new_n371_ & ~new_n370_ & new_n373_ & new_n349_ & new_n491_ & new_n493_;
  assign new_n491_ = new_n322_ & new_n288_ & new_n492_ & new_n326_ & new_n275_ & new_n284_ & ~new_n280_ & new_n293_;
  assign new_n492_ = (~DATAI_2_ | (new_n257_ & ~new_n258_)) & (new_n272_ | ~new_n257_ | new_n258_) & (~new_n260_ | ~new_n257_ | new_n258_) & (~DATAI_1_ | (new_n257_ & ~new_n258_)) & (~DATAI_0_ | (new_n257_ & ~new_n258_)) & (~IR_REG_0__SCAN_IN | ~new_n257_ | new_n258_);
  assign new_n493_ = new_n346_ & new_n343_ & new_n304_ & new_n308_ & new_n359_ & new_n342_ & new_n312_ & new_n316_;
  assign new_n494_ = (new_n495_ | ~new_n474_ | ~new_n499_) & ~new_n496_ & (~new_n498_ | ~new_n435_) & (new_n474_ | ~REG2_REG_28__SCAN_IN);
  assign new_n495_ = (~REG0_REG_29__SCAN_IN | new_n252_ | ~new_n255_) & (~REG1_REG_29__SCAN_IN | new_n252_ | new_n255_) & (~REG2_REG_29__SCAN_IN | ~new_n252_ | ~new_n255_) & (~new_n252_ | new_n255_ | ~new_n434_ | ~REG3_REG_28__SCAN_IN);
  assign new_n496_ = new_n497_ & (~new_n434_ | ~REG3_REG_28__SCAN_IN) & (new_n434_ | REG3_REG_28__SCAN_IN);
  assign new_n497_ = new_n485_ & new_n487_;
  assign new_n498_ = (IR_REG_20__SCAN_IN | (~new_n245_ & IR_REG_31__SCAN_IN)) & (~IR_REG_20__SCAN_IN | new_n245_ | ~IR_REG_31__SCAN_IN) & new_n474_ & (IR_REG_31__SCAN_IN ? ((new_n245_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN) | (IR_REG_21__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN))) : ~IR_REG_21__SCAN_IN) & (~IR_REG_22__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (new_n245_ & ~IR_REG_22__SCAN_IN & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN) | (IR_REG_22__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN)));
  assign new_n499_ = new_n257_ & new_n469_;
  assign new_n500_ = (IR_REG_20__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN))) & (~IR_REG_19__SCAN_IN ^ ((IR_REG_18__SCAN_IN & IR_REG_31__SCAN_IN) | (~new_n350_ & IR_REG_31__SCAN_IN))) & new_n474_ & (IR_REG_31__SCAN_IN ? ((~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN) | (IR_REG_21__SCAN_IN & (IR_REG_20__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN))) : ~IR_REG_21__SCAN_IN) & (~IR_REG_22__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_22__SCAN_IN & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN) | (IR_REG_22__SCAN_IN & (IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN)));
  assign new_n501_ = (~new_n524_ | (new_n474_ & (new_n518_ | ~new_n520_))) & (new_n502_ | ~new_n527_) & (~new_n522_ | (~new_n513_ & new_n474_));
  assign new_n502_ = new_n506_ & (~new_n503_ | new_n511_) & new_n507_ & (~new_n503_ | ~new_n512_);
  assign new_n503_ = new_n505_ ^ ((~new_n368_ & new_n370_) | ((~new_n368_ | new_n370_) & ~new_n373_ & ~new_n374_) | ((~new_n373_ | ~new_n374_) & (~new_n368_ | new_n370_) & ((~new_n349_ & ~new_n352_) | (~new_n504_ & (~new_n349_ | ~new_n352_)))));
  assign new_n504_ = new_n426_ & (~new_n420_ | (new_n418_ & (~new_n416_ | (~new_n421_ & (~new_n423_ | (new_n409_ & ~new_n422_))))));
  assign new_n505_ = new_n364_ ^ (new_n351_ | ~DATAI_21_);
  assign new_n506_ = (new_n368_ | ~new_n468_) & ((new_n441_ & ~new_n505_) | new_n470_ | (~new_n441_ & new_n505_));
  assign new_n507_ = (~new_n509_ | (new_n508_ & ~new_n371_) | (~new_n508_ & new_n371_)) & (~new_n371_ | ~new_n510_) & (new_n377_ | ~new_n499_);
  assign new_n508_ = ~new_n370_ & new_n373_ & new_n349_ & new_n491_ & new_n493_;
  assign new_n509_ = (IR_REG_31__SCAN_IN ? ((IR_REG_21__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN)) | (new_n245_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN)) : ~IR_REG_21__SCAN_IN) & (~IR_REG_22__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (new_n245_ & ~IR_REG_22__SCAN_IN & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN) | (IR_REG_22__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN))) & (IR_REG_20__SCAN_IN ^ (new_n245_ | ~IR_REG_31__SCAN_IN));
  assign new_n510_ = (IR_REG_31__SCAN_IN ? ((IR_REG_21__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN)) | (new_n245_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN)) : ~IR_REG_21__SCAN_IN) & (~IR_REG_22__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (new_n245_ & ~IR_REG_22__SCAN_IN & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN) | (IR_REG_22__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN))) & (IR_REG_20__SCAN_IN | (~new_n245_ & IR_REG_31__SCAN_IN)) & (~IR_REG_20__SCAN_IN | new_n245_ | ~IR_REG_31__SCAN_IN);
  assign new_n511_ = (new_n248_ | new_n249_ | (~new_n471_ & (IR_REG_21__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | ((~new_n245_ | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN) & (~IR_REG_21__SCAN_IN | (new_n245_ & ~IR_REG_20__SCAN_IN)))))) & ((~IR_REG_21__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & ((new_n245_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN) | (IR_REG_21__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN)))) | new_n248_ | new_n471_ | ~new_n249_);
  assign new_n512_ = new_n248_ & ~new_n471_ & new_n249_;
  assign new_n513_ = ((~new_n514_ & ~new_n516_) | new_n517_ | (new_n514_ & new_n516_)) & (((~new_n515_ | (~new_n377_ & ~new_n380_)) & (~new_n516_ | (new_n377_ & new_n380_))) | new_n470_ | (new_n516_ & new_n515_ & (new_n377_ | new_n380_))) & (new_n377_ | ~new_n468_) & (new_n516_ | new_n470_ | ~new_n377_ | ~new_n380_);
  assign new_n514_ = (~new_n377_ | new_n380_) & (new_n406_ | ~new_n424_ | (~new_n377_ & new_n380_));
  assign new_n515_ = (new_n364_ | new_n371_) & (~new_n441_ | (new_n364_ & new_n371_));
  assign new_n516_ = ~new_n382_ ^ new_n386_;
  assign new_n517_ = (((IR_REG_31__SCAN_IN ? ((~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN) | (IR_REG_21__SCAN_IN & (IR_REG_20__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN))) : ~IR_REG_21__SCAN_IN) & (~IR_REG_22__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_22__SCAN_IN & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN) | (IR_REG_22__SCAN_IN & (IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN)))) | ((~IR_REG_31__SCAN_IN | ((IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN) & (~IR_REG_21__SCAN_IN | (~IR_REG_20__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN)))) & (IR_REG_21__SCAN_IN | IR_REG_31__SCAN_IN) & ((IR_REG_22__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & (IR_REG_22__SCAN_IN | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN) & (~IR_REG_22__SCAN_IN | (~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN))))) | (~IR_REG_20__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN))) | (IR_REG_19__SCAN_IN ^ ((~new_n350_ & IR_REG_31__SCAN_IN) | (IR_REG_18__SCAN_IN & IR_REG_31__SCAN_IN)))) & ((~IR_REG_20__SCAN_IN & (~IR_REG_31__SCAN_IN | (new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN))) | (IR_REG_20__SCAN_IN & IR_REG_31__SCAN_IN & (~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN)) | ((~IR_REG_22__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_22__SCAN_IN & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN) | (IR_REG_22__SCAN_IN & (IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN)))) | (IR_REG_19__SCAN_IN ^ ((~new_n350_ & IR_REG_31__SCAN_IN) | (IR_REG_18__SCAN_IN & IR_REG_31__SCAN_IN)))) & ((IR_REG_19__SCAN_IN & ((~new_n350_ & IR_REG_31__SCAN_IN) | (IR_REG_18__SCAN_IN & IR_REG_31__SCAN_IN))) | (~IR_REG_19__SCAN_IN & (new_n350_ | ~IR_REG_31__SCAN_IN) & (~IR_REG_18__SCAN_IN | ~IR_REG_31__SCAN_IN)) | (IR_REG_31__SCAN_IN & ((~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN) | (IR_REG_21__SCAN_IN & (IR_REG_20__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN)))) | (~IR_REG_21__SCAN_IN & ~IR_REG_31__SCAN_IN) | (~IR_REG_20__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN))));
  assign new_n518_ = (new_n519_ | (~new_n373_ & ~new_n374_) | ((~new_n373_ | ~new_n374_) & ((~new_n349_ & ~new_n352_) | (~new_n504_ & (~new_n349_ | ~new_n352_))))) & ~new_n517_ & (~new_n519_ | ((new_n373_ | new_n374_) & ((new_n373_ & new_n374_) | ((new_n349_ | new_n352_) & (new_n504_ | (new_n349_ & new_n352_))))));
  assign new_n519_ = ~new_n368_ ^ new_n370_;
  assign new_n520_ = (new_n374_ | ~new_n468_) & ((new_n519_ & (~new_n373_ | new_n374_) & ((new_n521_ & (~new_n349_ | new_n352_)) | (~new_n349_ & new_n352_) | (~new_n373_ & new_n374_))) | new_n470_ | (~new_n519_ & ((new_n373_ & ~new_n374_) | ((~new_n521_ | (new_n349_ & ~new_n352_)) & (new_n349_ | ~new_n352_) & (new_n373_ | ~new_n374_)))));
  assign new_n521_ = new_n457_ & (~new_n455_ | (~new_n444_ & new_n453_));
  assign new_n522_ = new_n523_ & ((~new_n490_ & new_n386_) | ~new_n500_ | (new_n490_ & ~new_n386_));
  assign new_n523_ = (new_n396_ | ~new_n474_ | ~new_n499_) & (~new_n383_ | ~new_n497_) & (~new_n498_ | ~new_n386_) & (new_n474_ | ~REG2_REG_23__SCAN_IN);
  assign new_n524_ = ((new_n370_ & (~new_n373_ | ~new_n525_ | ~new_n349_)) | ~new_n500_ | (~new_n370_ & new_n373_ & new_n525_ & new_n349_)) & new_n526_ & (~new_n498_ | ~new_n370_);
  assign new_n525_ = new_n491_ & new_n493_;
  assign new_n526_ = (new_n364_ | ~new_n474_ | ~new_n499_) & (~new_n497_ | ~new_n369_) & (new_n474_ | ~REG2_REG_20__SCAN_IN);
  assign new_n527_ = new_n475_ & ~new_n529_ & new_n485_ & ~new_n528_ & ~new_n487_ & ~new_n488_;
  assign new_n528_ = ~new_n480_ & (~new_n476_ | new_n477_ | ~B_REG_SCAN_IN) & ~new_n478_ & (~new_n477_ | B_REG_SCAN_IN);
  assign new_n529_ = (~new_n476_ | ~new_n478_) & (D_REG_1__SCAN_IN | (new_n476_ & ~new_n477_ & B_REG_SCAN_IN) | new_n478_ | (new_n477_ & ~B_REG_SCAN_IN));
  assign new_n530_ = ~new_n531_ & ~new_n539_ & new_n647_ & new_n542_ & new_n564_ & ~new_n652_ & (~new_n649_ | ~new_n618_);
  assign new_n531_ = ((~new_n533_ & (new_n391_ | new_n393_) & (~new_n391_ | ~new_n393_)) | new_n538_ | (new_n533_ & (new_n391_ ^ ~new_n393_))) & new_n535_ & ((new_n532_ & (new_n391_ ^ ~new_n393_)) | new_n470_ | (~new_n532_ & (new_n391_ | new_n393_) & (~new_n391_ | ~new_n393_)));
  assign new_n532_ = ~new_n467_ & (~new_n464_ | (new_n462_ & (~new_n441_ | ~new_n461_)));
  assign new_n533_ = ~new_n429_ & (~new_n534_ | (new_n428_ & (new_n405_ | ((~new_n377_ | new_n380_) & (new_n406_ | ~new_n424_ | (~new_n377_ & new_n380_))))));
  assign new_n534_ = (new_n394_ | ~new_n395_) & (new_n396_ | ~new_n399_);
  assign new_n535_ = new_n536_ & ((~new_n393_ & ~new_n395_ & ~new_n399_ & new_n490_ & ~new_n386_) | ~new_n509_ | (new_n393_ & (new_n395_ | new_n399_ | ~new_n490_ | new_n386_)));
  assign new_n536_ = (new_n431_ | ~new_n499_) & (new_n394_ | ~new_n468_) & new_n537_ & (~new_n393_ | ~new_n510_);
  assign new_n537_ = ~new_n475_ & ~new_n529_ & new_n485_ & ~new_n528_ & ~new_n487_ & ~new_n488_;
  assign new_n538_ = (((IR_REG_31__SCAN_IN ? ((~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN) | (IR_REG_21__SCAN_IN & (IR_REG_20__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN))) : ~IR_REG_21__SCAN_IN) & (~IR_REG_22__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_22__SCAN_IN & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN) | (IR_REG_22__SCAN_IN & (IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN)))) | ((~IR_REG_31__SCAN_IN | ((IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN) & (~IR_REG_21__SCAN_IN | (~IR_REG_20__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN)))) & (IR_REG_21__SCAN_IN | IR_REG_31__SCAN_IN) & ((IR_REG_22__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & (IR_REG_22__SCAN_IN | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN) & (~IR_REG_22__SCAN_IN | (~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN))))) | (~IR_REG_20__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN))) | (IR_REG_19__SCAN_IN ^ ((~new_n350_ & IR_REG_31__SCAN_IN) | (IR_REG_18__SCAN_IN & IR_REG_31__SCAN_IN)))) & ((~IR_REG_20__SCAN_IN & (~IR_REG_31__SCAN_IN | (new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN))) | (IR_REG_20__SCAN_IN & IR_REG_31__SCAN_IN & (~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN)) | ((~IR_REG_22__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_22__SCAN_IN & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN) | (IR_REG_22__SCAN_IN & (IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN)))) | (IR_REG_19__SCAN_IN ^ ((~new_n350_ & IR_REG_31__SCAN_IN) | (IR_REG_18__SCAN_IN & IR_REG_31__SCAN_IN)))) & ((IR_REG_19__SCAN_IN & ((~new_n350_ & IR_REG_31__SCAN_IN) | (IR_REG_18__SCAN_IN & IR_REG_31__SCAN_IN))) | (~IR_REG_19__SCAN_IN & (new_n350_ | ~IR_REG_31__SCAN_IN) & (~IR_REG_18__SCAN_IN | ~IR_REG_31__SCAN_IN)) | (IR_REG_22__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & (IR_REG_22__SCAN_IN | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN | ~new_n350_ | IR_REG_18__SCAN_IN | IR_REG_19__SCAN_IN) & (~IR_REG_22__SCAN_IN | (~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN & new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN))) | (~IR_REG_20__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (new_n350_ & ~IR_REG_18__SCAN_IN & ~IR_REG_19__SCAN_IN))));
  assign new_n539_ = new_n474_ & (~new_n506_ | (new_n503_ & ~new_n511_) | ~new_n540_ | ((new_n515_ | ~new_n541_) & ~new_n470_ & (~new_n515_ | new_n541_)));
  assign new_n540_ = (new_n364_ | ~new_n468_) & (new_n436_ | (new_n541_ ^ (new_n406_ | ~new_n424_)));
  assign new_n541_ = new_n377_ ^ new_n380_;
  assign new_n542_ = ((~new_n543_ & new_n563_) | ~new_n555_ | (new_n543_ & ~new_n563_)) & ~new_n544_ & (~new_n560_ | (~new_n557_ & new_n474_));
  assign new_n543_ = (new_n356_ | new_n360_) & ((new_n356_ & new_n360_) | (~new_n236_ & new_n330_));
  assign new_n544_ = new_n547_ & (~new_n555_ | (~new_n556_ ^ (new_n333_ | (~new_n545_ & ~new_n301_))));
  assign new_n545_ = ~new_n546_ & (new_n319_ | (~new_n296_ & (~new_n276_ | (~new_n324_ & (new_n237_ | ~new_n328_))))) & (new_n329_ | (new_n319_ & ~new_n296_ & (~new_n276_ | (~new_n324_ & (new_n237_ | ~new_n328_)))));
  assign new_n546_ = ((new_n239_ & ~new_n302_) | (new_n250_ & ~new_n304_)) & (new_n269_ ^ ((new_n250_ & ~new_n302_) | (new_n262_ & ~new_n304_)));
  assign new_n547_ = (new_n548_ | (REG3_REG_12__SCAN_IN & new_n307_ & REG3_REG_11__SCAN_IN) | (~REG3_REG_12__SCAN_IN & (~new_n307_ | ~REG3_REG_11__SCAN_IN))) & (~new_n553_ | new_n312_) & ~new_n554_ & (STATE_REG_SCAN_IN | ~REG3_REG_12__SCAN_IN);
  assign new_n548_ = ~new_n549_ & (new_n550_ | ~new_n552_);
  assign new_n549_ = STATE_REG_SCAN_IN & ((~new_n550_ & new_n510_) | (~new_n550_ & ~new_n551_) | new_n488_ | new_n240_ | new_n486_);
  assign new_n550_ = (new_n477_ | ~new_n478_) & (D_REG_0__SCAN_IN | (new_n476_ & ~new_n477_ & B_REG_SCAN_IN) | new_n478_ | (new_n477_ & ~B_REG_SCAN_IN)) & (new_n480_ | (new_n476_ & ~new_n477_ & B_REG_SCAN_IN) | new_n478_ | (new_n477_ & ~B_REG_SCAN_IN)) & (~new_n476_ | ~new_n478_) & (D_REG_1__SCAN_IN | (new_n476_ & ~new_n477_ & B_REG_SCAN_IN) | new_n478_ | (new_n477_ & ~B_REG_SCAN_IN));
  assign new_n551_ = (((IR_REG_22__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & (~new_n245_ | IR_REG_22__SCAN_IN | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN) & (~IR_REG_22__SCAN_IN | (new_n245_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN)))) ^ (IR_REG_31__SCAN_IN ? ((new_n245_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN) | (IR_REG_21__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN))) : ~IR_REG_21__SCAN_IN)) & (new_n248_ | (IR_REG_22__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & (~new_n245_ | IR_REG_22__SCAN_IN | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN) & (~IR_REG_22__SCAN_IN | (new_n245_ & ~IR_REG_20__SCAN_IN & ~IR_REG_21__SCAN_IN))) | (~IR_REG_20__SCAN_IN ^ (new_n245_ | ~IR_REG_31__SCAN_IN)));
  assign new_n552_ = new_n469_ & ~new_n248_ & ~new_n471_ & STATE_REG_SCAN_IN & ~new_n240_ & ~new_n486_;
  assign new_n553_ = new_n485_ & (new_n487_ | (new_n550_ & new_n510_));
  assign new_n554_ = new_n552_ & ((~new_n306_ & new_n550_ & ~new_n257_) | (~new_n314_ & new_n550_ & new_n257_));
  assign new_n555_ = new_n550_ & new_n485_ & ~new_n551_;
  assign new_n556_ = ((~new_n239_ | new_n311_) & (~new_n250_ | new_n312_)) ^ (~new_n269_ ^ ((new_n250_ & ~new_n311_) | (new_n262_ & ~new_n312_)));
  assign new_n557_ = (new_n511_ | (new_n504_ & ~new_n558_) | (~new_n504_ & new_n558_)) & ~new_n559_ & ((new_n521_ & new_n558_) | new_n470_ | (~new_n521_ & ~new_n558_));
  assign new_n558_ = new_n349_ ^ new_n352_;
  assign new_n559_ = ~new_n336_ & new_n468_;
  assign new_n560_ = (~new_n473_ | (~new_n504_ & (new_n349_ | new_n352_) & (~new_n349_ | ~new_n352_)) | (new_n504_ & (new_n349_ ^ ~new_n352_))) & new_n561_ & (~new_n500_ | (new_n525_ & new_n349_) | (~new_n525_ & ~new_n349_));
  assign new_n561_ = (new_n562_ | ~new_n474_) & (new_n474_ | ~REG2_REG_18__SCAN_IN) & (~new_n497_ | (new_n353_ & REG3_REG_18__SCAN_IN) | (~new_n353_ & ~REG3_REG_18__SCAN_IN));
  assign new_n562_ = (new_n374_ | ~new_n499_) & (new_n349_ | ~new_n510_);
  assign new_n563_ = ((~new_n239_ | new_n340_) & (~new_n250_ | new_n342_)) ^ (~new_n269_ ^ ((new_n250_ & ~new_n340_) | (new_n262_ & ~new_n342_)));
  assign new_n564_ = ~new_n565_ & (~new_n567_ | ~new_n618_) & new_n582_ & (~new_n644_ | (new_n555_ & (~new_n643_ ^ ~new_n646_)));
  assign new_n565_ = (new_n511_ | (new_n504_ & ~new_n558_) | (~new_n504_ & new_n558_)) & ~new_n559_ & ((new_n521_ & new_n558_) | new_n470_ | (~new_n521_ & ~new_n558_)) & new_n566_ & (~new_n512_ | (new_n504_ & ~new_n558_) | (~new_n504_ & new_n558_));
  assign new_n566_ = new_n562_ & new_n537_ & (~new_n509_ | (new_n525_ & new_n349_) | (~new_n525_ & ~new_n349_));
  assign new_n567_ = ~new_n258_ & (new_n568_ ^ (~new_n344_ ^ ~REG1_REG_17__SCAN_IN));
  assign new_n568_ = (new_n581_ | REG1_REG_16__SCAN_IN) & ((new_n581_ & REG1_REG_16__SCAN_IN) | ((new_n580_ | REG1_REG_15__SCAN_IN) & ((new_n580_ & REG1_REG_15__SCAN_IN) | (~new_n569_ & (~new_n571_ | REG1_REG_14__SCAN_IN)))));
  assign new_n569_ = ~new_n570_ & ((new_n579_ & ~REG1_REG_13__SCAN_IN) | ((new_n579_ | ~REG1_REG_13__SCAN_IN) & ((~new_n313_ & ~REG1_REG_12__SCAN_IN) | ((~new_n572_ | (~new_n309_ & ~REG1_REG_11__SCAN_IN)) & (~new_n309_ | ~REG1_REG_11__SCAN_IN) & (~new_n313_ | ~REG1_REG_12__SCAN_IN)))));
  assign new_n570_ = ~new_n571_ & REG1_REG_14__SCAN_IN;
  assign new_n571_ = IR_REG_14__SCAN_IN ^ (new_n317_ | ~IR_REG_31__SCAN_IN);
  assign new_n572_ = (~new_n305_ | REG1_REG_10__SCAN_IN) & ((~new_n305_ & REG1_REG_10__SCAN_IN) | ((~new_n323_ | REG1_REG_9__SCAN_IN) & ((~new_n323_ & REG1_REG_9__SCAN_IN) | ((~new_n294_ | REG1_REG_8__SCAN_IN) & (new_n573_ | (~new_n294_ & REG1_REG_8__SCAN_IN))))));
  assign new_n573_ = (new_n281_ | REG1_REG_7__SCAN_IN) & (new_n574_ | (~new_n285_ & REG1_REG_6__SCAN_IN) | (new_n281_ & REG1_REG_7__SCAN_IN));
  assign new_n574_ = (~new_n285_ | REG1_REG_6__SCAN_IN) & ((new_n289_ & REG1_REG_5__SCAN_IN) | ((~new_n577_ | (~new_n575_ & new_n576_)) & ~new_n578_ & (new_n289_ | REG1_REG_5__SCAN_IN)));
  assign new_n575_ = (~REG1_REG_2__SCAN_IN | ((~IR_REG_2__SCAN_IN | IR_REG_31__SCAN_IN) & (~IR_REG_31__SCAN_IN | (~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN) | (IR_REG_2__SCAN_IN & (IR_REG_0__SCAN_IN | IR_REG_1__SCAN_IN))))) & ((~REG1_REG_1__SCAN_IN & (~IR_REG_1__SCAN_IN ^ (IR_REG_0__SCAN_IN & IR_REG_31__SCAN_IN))) | ((~IR_REG_0__SCAN_IN | ~REG1_REG_0__SCAN_IN) & (~REG1_REG_1__SCAN_IN | (IR_REG_1__SCAN_IN & IR_REG_0__SCAN_IN & IR_REG_31__SCAN_IN) | (~IR_REG_1__SCAN_IN & (~IR_REG_0__SCAN_IN | ~IR_REG_31__SCAN_IN)))));
  assign new_n576_ = (REG1_REG_2__SCAN_IN | (IR_REG_2__SCAN_IN & ~IR_REG_31__SCAN_IN) | ((~IR_REG_2__SCAN_IN | (~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN)) & IR_REG_31__SCAN_IN & (IR_REG_2__SCAN_IN | IR_REG_0__SCAN_IN | IR_REG_1__SCAN_IN))) & (REG1_REG_3__SCAN_IN | (~IR_REG_3__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN))));
  assign new_n577_ = (~REG1_REG_3__SCAN_IN | (~IR_REG_3__SCAN_IN & (~IR_REG_31__SCAN_IN | (~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN))) | (IR_REG_3__SCAN_IN & IR_REG_31__SCAN_IN & (IR_REG_2__SCAN_IN | IR_REG_0__SCAN_IN | IR_REG_1__SCAN_IN))) & (~REG1_REG_4__SCAN_IN | (IR_REG_4__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_3__SCAN_IN & ~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN))));
  assign new_n578_ = ~REG1_REG_4__SCAN_IN & (~IR_REG_4__SCAN_IN | (IR_REG_31__SCAN_IN & (IR_REG_3__SCAN_IN | IR_REG_2__SCAN_IN | IR_REG_0__SCAN_IN | IR_REG_1__SCAN_IN))) & (IR_REG_4__SCAN_IN | ~IR_REG_31__SCAN_IN | (~IR_REG_3__SCAN_IN & ~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN));
  assign new_n579_ = (~IR_REG_13__SCAN_IN | IR_REG_31__SCAN_IN) & ((IR_REG_13__SCAN_IN & (~new_n318_ | IR_REG_12__SCAN_IN)) | new_n317_ | ~IR_REG_31__SCAN_IN);
  assign new_n580_ = (IR_REG_15__SCAN_IN | (IR_REG_31__SCAN_IN & (~new_n317_ | IR_REG_14__SCAN_IN))) & (~IR_REG_15__SCAN_IN | ~IR_REG_31__SCAN_IN | (new_n317_ & ~IR_REG_14__SCAN_IN));
  assign new_n581_ = IR_REG_16__SCAN_IN ^ ((IR_REG_15__SCAN_IN & IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & (~new_n317_ | IR_REG_14__SCAN_IN)));
  assign new_n582_ = ~new_n583_ & ~new_n589_ & new_n632_ & new_n626_ & new_n624_ & new_n623_ & ~new_n590_ & new_n594_;
  assign new_n583_ = new_n537_ & (((new_n409_ | new_n588_) & ~new_n538_ & (~new_n409_ | ~new_n588_)) | ~new_n586_ | ((new_n588_ | new_n584_ | ~new_n585_) & ~new_n470_ & (~new_n588_ | (~new_n584_ & new_n585_))));
  assign new_n584_ = new_n448_ & ~new_n445_ & new_n446_;
  assign new_n585_ = new_n450_ & (~new_n447_ | new_n449_);
  assign new_n586_ = ((~new_n587_ & ~new_n322_) | ~new_n509_ | (new_n587_ & new_n322_)) & (new_n302_ | ~new_n499_) & (new_n291_ | ~new_n468_) & (new_n322_ | ~new_n510_);
  assign new_n587_ = new_n288_ & new_n492_ & new_n326_ & new_n275_ & new_n284_ & ~new_n280_ & new_n293_;
  assign new_n588_ = ~new_n320_ ^ new_n322_;
  assign new_n589_ = new_n552_ & ((~new_n433_ & new_n550_ & new_n257_) | (new_n432_ & ~new_n550_) | (~new_n391_ & new_n550_ & ~new_n257_));
  assign new_n590_ = new_n527_ & ((~new_n470_ & (new_n593_ ^ (~new_n270_ ^ ~new_n271_))) | ~new_n591_ | ((~new_n411_ | (new_n270_ ^ ~new_n271_)) & ~new_n538_ & (new_n411_ | (new_n270_ & ~new_n271_) | (~new_n270_ & new_n271_))));
  assign new_n591_ = new_n592_ & ((~new_n271_ & (~new_n256_ | ~new_n264_)) | ~new_n509_ | (new_n271_ & new_n256_ & new_n264_));
  assign new_n592_ = (new_n251_ | ~new_n468_) & (new_n274_ | ~new_n499_) & (new_n271_ | ~new_n510_);
  assign new_n593_ = (~new_n256_ | (new_n251_ & ~new_n264_ & new_n265_)) & (new_n251_ | (~new_n264_ & new_n265_));
  assign new_n594_ = new_n619_ & (new_n548_ | ~REG3_REG_0__SCAN_IN) & new_n595_ & new_n613_ & (~new_n380_ | (~new_n498_ & ~new_n553_));
  assign new_n595_ = ~new_n598_ & new_n609_ & new_n599_ & (~new_n597_ | new_n612_) & (~new_n596_ | (~ADDR_REG_17__SCAN_IN & ~ADDR_REG_1__SCAN_IN));
  assign new_n596_ = STATE_REG_SCAN_IN & (~new_n240_ | new_n486_) & ((new_n240_ & ~new_n486_) | new_n351_ | (~new_n486_ & new_n469_));
  assign new_n597_ = STATE_REG_SCAN_IN & ~new_n240_ & ~new_n486_ & (~new_n240_ | new_n486_) & ~new_n351_ & (new_n486_ | ~new_n469_);
  assign new_n598_ = (REG2_REG_21__SCAN_IN | REG2_REG_22__SCAN_IN) & (~new_n485_ | (~new_n487_ & (~new_n479_ | new_n475_ | new_n488_)));
  assign new_n599_ = (~new_n485_ | ((~new_n476_ | new_n477_ | ~B_REG_SCAN_IN) & ~new_n478_ & (~new_n477_ | B_REG_SCAN_IN)) | new_n477_ | (new_n476_ & ~new_n478_)) & (new_n608_ | (new_n485_ & ((new_n476_ & ~new_n477_ & B_REG_SCAN_IN) | new_n478_ | (new_n477_ & ~B_REG_SCAN_IN)))) & new_n600_ & new_n605_ & (~new_n485_ | ((~new_n476_ | new_n477_ | ~B_REG_SCAN_IN) & ~new_n478_ & (~new_n477_ | B_REG_SCAN_IN)));
  assign new_n600_ = new_n602_ & ((DATAI_30_ & ~STATE_REG_SCAN_IN) | (IR_REG_30__SCAN_IN & STATE_REG_SCAN_IN & ~IR_REG_31__SCAN_IN) | (STATE_REG_SCAN_IN & IR_REG_31__SCAN_IN & (IR_REG_30__SCAN_IN | ~new_n601_ | ~new_n254_) & (~IR_REG_30__SCAN_IN | (new_n601_ & new_n254_))));
  assign new_n601_ = new_n253_ & new_n243_ & new_n244_ & new_n241_ & new_n242_;
  assign new_n602_ = ((DATAI_7_ & ~STATE_REG_SCAN_IN) | (IR_REG_7__SCAN_IN & STATE_REG_SCAN_IN & ~IR_REG_31__SCAN_IN) | (STATE_REG_SCAN_IN & IR_REG_31__SCAN_IN & (new_n241_ | ~IR_REG_7__SCAN_IN) & (~new_n241_ | IR_REG_7__SCAN_IN))) & (new_n604_ | STATE_REG_SCAN_IN) & D_REG_14__SCAN_IN & (new_n603_ | ~STATE_REG_SCAN_IN | IR_REG_31__SCAN_IN);
  assign new_n603_ = ~IR_REG_24__SCAN_IN & ~IR_REG_27__SCAN_IN;
  assign new_n604_ = ~REG3_REG_27__SCAN_IN & ~REG3_REG_1__SCAN_IN & ~DATAI_27_ & ~DATAI_24_ & ~REG3_REG_17__SCAN_IN & ~REG3_REG_0__SCAN_IN & ~REG3_REG_15__SCAN_IN & ~REG3_REG_22__SCAN_IN;
  assign new_n605_ = ~new_n606_ & ((STATE_REG_SCAN_IN & IR_REG_31__SCAN_IN & (~new_n245_ | IR_REG_20__SCAN_IN | IR_REG_21__SCAN_IN) & (~IR_REG_21__SCAN_IN | (new_n245_ & ~IR_REG_20__SCAN_IN))) | (DATAI_21_ & ~STATE_REG_SCAN_IN) | (IR_REG_21__SCAN_IN & STATE_REG_SCAN_IN & ~IR_REG_31__SCAN_IN)) & (new_n607_ | ~STATE_REG_SCAN_IN | ~IR_REG_31__SCAN_IN);
  assign new_n606_ = (~STATE_REG_SCAN_IN | ~IR_REG_31__SCAN_IN | (~IR_REG_11__SCAN_IN & ~IR_REG_10__SCAN_IN & ~IR_REG_9__SCAN_IN & new_n295_ & ~IR_REG_8__SCAN_IN) | (IR_REG_11__SCAN_IN & (IR_REG_10__SCAN_IN | IR_REG_9__SCAN_IN | ~new_n295_ | IR_REG_8__SCAN_IN))) & (~DATAI_11_ | STATE_REG_SCAN_IN) & (~IR_REG_11__SCAN_IN | ~STATE_REG_SCAN_IN | IR_REG_31__SCAN_IN);
  assign new_n607_ = ((new_n243_ & new_n244_ & new_n241_ & new_n242_ & new_n259_ & ~IR_REG_24__SCAN_IN & ~IR_REG_27__SCAN_IN) | (IR_REG_27__SCAN_IN & (~new_n259_ | IR_REG_24__SCAN_IN | ~new_n243_ | ~new_n244_ | ~new_n241_ | ~new_n242_))) & (IR_REG_24__SCAN_IN ^ (new_n243_ & new_n244_ & new_n241_ & new_n242_));
  assign new_n608_ = ~D_REG_4__SCAN_IN & ~D_REG_8__SCAN_IN & ~D_REG_27__SCAN_IN & ~D_REG_31__SCAN_IN & D_REG_0__SCAN_IN & ~D_REG_18__SCAN_IN;
  assign new_n609_ = (new_n610_ | (new_n475_ & ~new_n529_ & new_n485_ & ~new_n528_ & ~new_n487_ & ~new_n488_)) & (new_n611_ | (~new_n475_ & ~new_n529_ & new_n485_ & ~new_n528_ & ~new_n487_ & ~new_n488_));
  assign new_n610_ = ~REG1_REG_21__SCAN_IN & ~REG1_REG_2__SCAN_IN & REG1_REG_5__SCAN_IN;
  assign new_n611_ = ~REG0_REG_9__SCAN_IN & REG0_REG_18__SCAN_IN & REG0_REG_29__SCAN_IN & REG0_REG_26__SCAN_IN & ~REG0_REG_27__SCAN_IN;
  assign new_n612_ = (new_n257_ | ~new_n258_ | (~REG2_REG_1__SCAN_IN & (~new_n260_ ^ (IR_REG_0__SCAN_IN & REG2_REG_0__SCAN_IN))) | (REG2_REG_1__SCAN_IN & (~new_n260_ | ~IR_REG_0__SCAN_IN | ~REG2_REG_0__SCAN_IN) & (new_n260_ | (IR_REG_0__SCAN_IN & REG2_REG_0__SCAN_IN)))) & (~new_n257_ | ~new_n260_) & (new_n258_ | ((~IR_REG_0__SCAN_IN | ~REG1_REG_0__SCAN_IN) & (~new_n260_ ^ REG1_REG_1__SCAN_IN)) | (IR_REG_0__SCAN_IN & REG1_REG_0__SCAN_IN & (~new_n260_ | ~REG1_REG_1__SCAN_IN) & (new_n260_ | REG1_REG_1__SCAN_IN)));
  assign new_n613_ = ~new_n614_ & ~new_n615_ & new_n617_;
  assign new_n614_ = (~new_n264_ | ~new_n342_ | new_n437_) & new_n485_ & (new_n487_ | (new_n550_ & new_n510_));
  assign new_n615_ = (new_n278_ | new_n302_ | ~new_n616_) & (new_n616_ | ~DATAO_REG_7__SCAN_IN | ~DATAO_REG_10__SCAN_IN | ~DATAO_REG_26__SCAN_IN | DATAO_REG_21__SCAN_IN | DATAO_REG_22__SCAN_IN);
  assign new_n616_ = STATE_REG_SCAN_IN & new_n240_ & ~new_n486_;
  assign new_n617_ = (~new_n550_ | ~new_n257_ | new_n251_ | ~new_n552_) & (~new_n618_ | (new_n612_ & (~new_n257_ | ~new_n344_)));
  assign new_n618_ = new_n486_ & STATE_REG_SCAN_IN & (((~new_n240_ | new_n486_) & (~new_n257_ | new_n258_) & (new_n486_ | ~new_n469_)) | ~STATE_REG_SCAN_IN | (new_n240_ & ~new_n486_));
  assign new_n619_ = ~new_n620_ & (~new_n549_ | ~new_n341_) & (new_n621_ | new_n267_ | ~new_n555_) & ~new_n622_ & (~new_n549_ | ~new_n378_);
  assign new_n620_ = (new_n616_ | ~DATAO_REG_19__SCAN_IN) & (~new_n379_ | (new_n365_ & new_n378_) | ~new_n367_ | (new_n365_ & new_n366_) | new_n374_ | ~new_n616_);
  assign new_n621_ = (~new_n250_ | new_n265_) & (~new_n262_ | new_n264_) & (~new_n240_ | ~REG1_REG_0__SCAN_IN) & (~new_n240_ | ~IR_REG_0__SCAN_IN) & (~new_n250_ | new_n264_) & (~new_n239_ | new_n265_);
  assign new_n622_ = new_n552_ & ((~new_n345_ & new_n550_ & new_n257_) | (~new_n550_ & new_n341_) | (~new_n357_ & new_n550_ & ~new_n257_));
  assign new_n623_ = (~new_n432_ | ~new_n549_) & (~new_n552_ | ((new_n382_ | ~new_n550_ | ~new_n257_) & (~new_n378_ | new_n550_) & (new_n364_ | ~new_n550_ | new_n257_)));
  assign new_n624_ = (~new_n391_ | ~new_n616_) & (~new_n474_ | (new_n625_ & (~new_n499_ | (new_n382_ & new_n377_))));
  assign new_n625_ = (~new_n371_ | ~new_n510_) & (~new_n487_ | (~new_n366_ & ~new_n378_));
  assign new_n626_ = (~new_n500_ | (~new_n508_ & new_n371_) | (new_n508_ & ~new_n371_)) & ((~new_n627_ & ~new_n470_) | new_n628_ | ~new_n630_);
  assign new_n627_ = ((new_n445_ | ~new_n446_) & (new_n325_ | ~new_n326_)) ^ (~new_n287_ ^ new_n288_);
  assign new_n628_ = ((~new_n287_ & ~new_n288_) | (new_n287_ & new_n288_) | (new_n325_ & new_n326_) | (~new_n629_ & (new_n274_ | new_n275_) & (new_n325_ | new_n326_))) & ~new_n538_ & ((~new_n287_ ^ ~new_n288_) | ((~new_n325_ | ~new_n326_) & (new_n629_ | (~new_n274_ & ~new_n275_) | (~new_n325_ & ~new_n326_))));
  assign new_n629_ = (~new_n270_ | ~new_n271_) & (~new_n274_ | ~new_n275_) & ((~new_n270_ & ~new_n271_) | ((~new_n251_ | ~new_n256_) & ((~new_n264_ & ~new_n265_) | (~new_n251_ & ~new_n256_))));
  assign new_n630_ = new_n527_ & new_n631_ & ((~new_n288_ & (~new_n492_ | ~new_n326_ | ~new_n275_)) | ~new_n509_ | (new_n288_ & new_n492_ & new_n326_ & new_n275_));
  assign new_n631_ = (new_n325_ | ~new_n468_) & (new_n283_ | ~new_n499_) & (new_n288_ | ~new_n510_);
  assign new_n632_ = ((~new_n633_ & new_n380_) | ~new_n500_ | (new_n633_ & ~new_n380_)) & (new_n634_ | (new_n596_ & ADDR_REG_11__SCAN_IN) | (~STATE_REG_SCAN_IN & REG3_REG_11__SCAN_IN));
  assign new_n633_ = ~new_n371_ & ~new_n370_ & new_n373_ & new_n349_ & new_n491_ & new_n493_;
  assign new_n634_ = (new_n597_ | new_n618_) & (new_n635_ | (new_n257_ & new_n309_) | ((~new_n572_ | (~new_n309_ & ~REG1_REG_11__SCAN_IN) | (new_n309_ & REG1_REG_11__SCAN_IN)) & ~new_n258_ & (new_n572_ | (~new_n309_ ^ ~REG1_REG_11__SCAN_IN))));
  assign new_n635_ = ((new_n309_ & REG2_REG_11__SCAN_IN) | (~new_n309_ & ~REG2_REG_11__SCAN_IN) | ((new_n305_ | ~REG2_REG_10__SCAN_IN) & (new_n636_ | (new_n305_ & ~REG2_REG_10__SCAN_IN)))) & new_n642_ & ((new_n309_ ^ REG2_REG_11__SCAN_IN) | (~new_n305_ & REG2_REG_10__SCAN_IN) | (~new_n636_ & (~new_n305_ | REG2_REG_10__SCAN_IN)));
  assign new_n636_ = (new_n323_ | ~REG2_REG_9__SCAN_IN) & ((new_n323_ & ~REG2_REG_9__SCAN_IN) | ((new_n294_ | ~REG2_REG_8__SCAN_IN) & ((new_n294_ & ~REG2_REG_8__SCAN_IN) | ((~new_n281_ | ~REG2_REG_7__SCAN_IN) & (new_n637_ | (~new_n281_ & ~REG2_REG_7__SCAN_IN))))));
  assign new_n637_ = (new_n285_ | ~REG2_REG_6__SCAN_IN) & ((new_n285_ & ~REG2_REG_6__SCAN_IN) | ((~new_n289_ | ~REG2_REG_5__SCAN_IN) & ((~new_n289_ & ~REG2_REG_5__SCAN_IN) | (~new_n638_ & (~new_n641_ | (~new_n639_ & new_n640_))))));
  assign new_n638_ = REG2_REG_4__SCAN_IN & (~IR_REG_4__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_3__SCAN_IN & ~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN)));
  assign new_n639_ = (REG2_REG_2__SCAN_IN | (IR_REG_2__SCAN_IN & ~IR_REG_31__SCAN_IN) | (IR_REG_31__SCAN_IN & (IR_REG_2__SCAN_IN | IR_REG_0__SCAN_IN | IR_REG_1__SCAN_IN) & (~IR_REG_2__SCAN_IN | (~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN)))) & (REG2_REG_1__SCAN_IN | (IR_REG_0__SCAN_IN & REG2_REG_0__SCAN_IN & (~IR_REG_1__SCAN_IN | ~IR_REG_0__SCAN_IN | ~IR_REG_31__SCAN_IN) & (IR_REG_1__SCAN_IN | (IR_REG_0__SCAN_IN & IR_REG_31__SCAN_IN)))) & ((IR_REG_0__SCAN_IN & REG2_REG_0__SCAN_IN) | (IR_REG_1__SCAN_IN ^ (IR_REG_0__SCAN_IN & IR_REG_31__SCAN_IN)));
  assign new_n640_ = (~REG2_REG_3__SCAN_IN | (~IR_REG_3__SCAN_IN & (~IR_REG_31__SCAN_IN | (~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN))) | (IR_REG_3__SCAN_IN & IR_REG_31__SCAN_IN & (IR_REG_2__SCAN_IN | IR_REG_0__SCAN_IN | IR_REG_1__SCAN_IN))) & (~REG2_REG_2__SCAN_IN | ((~IR_REG_2__SCAN_IN | IR_REG_31__SCAN_IN) & ((IR_REG_2__SCAN_IN & (IR_REG_0__SCAN_IN | IR_REG_1__SCAN_IN)) | ~IR_REG_31__SCAN_IN | (~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN))));
  assign new_n641_ = (REG2_REG_4__SCAN_IN | (IR_REG_4__SCAN_IN & (~IR_REG_31__SCAN_IN | (~IR_REG_3__SCAN_IN & ~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN))) | (~IR_REG_4__SCAN_IN & IR_REG_31__SCAN_IN & (IR_REG_3__SCAN_IN | IR_REG_2__SCAN_IN | IR_REG_0__SCAN_IN | IR_REG_1__SCAN_IN))) & (REG2_REG_3__SCAN_IN | (~IR_REG_3__SCAN_IN ^ (~IR_REG_31__SCAN_IN | (~IR_REG_2__SCAN_IN & ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN))));
  assign new_n642_ = ~new_n257_ & new_n258_;
  assign new_n643_ = ~new_n282_ & (new_n297_ | new_n298_ | (~new_n286_ & (new_n324_ | (~new_n237_ & new_n328_))));
  assign new_n644_ = (new_n548_ | (~REG3_REG_7__SCAN_IN & (~new_n279_ | ~REG3_REG_6__SCAN_IN)) | (new_n279_ & REG3_REG_7__SCAN_IN & REG3_REG_6__SCAN_IN)) & (~new_n553_ | ~new_n280_) & ~new_n645_ & (STATE_REG_SCAN_IN | ~REG3_REG_7__SCAN_IN);
  assign new_n645_ = new_n552_ & ((~new_n283_ & new_n550_ & ~new_n257_) | (~new_n291_ & new_n550_ & new_n257_));
  assign new_n646_ = (~new_n269_ ^ ((new_n250_ & ~new_n278_) | (new_n262_ & new_n280_))) ^ ((~new_n239_ | new_n278_) & (~new_n250_ | ~new_n280_));
  assign new_n647_ = ~new_n648_ & (~new_n473_ | (~new_n503_ & (~new_n541_ | (~new_n406_ & new_n424_)) & (new_n541_ | new_n406_ | ~new_n424_)));
  assign new_n648_ = new_n597_ & (new_n649_ | (new_n257_ & new_n344_) | (~new_n258_ & (new_n568_ ^ (~new_n344_ ^ ~REG1_REG_17__SCAN_IN))));
  assign new_n649_ = (new_n344_ | (REG2_REG_17__SCAN_IN & ((~new_n581_ & ~REG2_REG_16__SCAN_IN) | (new_n650_ & (~new_n581_ | ~REG2_REG_16__SCAN_IN)))) | (~REG2_REG_17__SCAN_IN & (new_n581_ | REG2_REG_16__SCAN_IN) & (~new_n650_ | (new_n581_ & REG2_REG_16__SCAN_IN)))) & new_n642_ & (~new_n344_ | (REG2_REG_17__SCAN_IN ^ ((~new_n581_ & ~REG2_REG_16__SCAN_IN) | (new_n650_ & (~new_n581_ | ~REG2_REG_16__SCAN_IN)))));
  assign new_n650_ = (~new_n580_ | ~REG2_REG_15__SCAN_IN) & ((~new_n580_ & ~REG2_REG_15__SCAN_IN) | ((new_n571_ | ~REG2_REG_14__SCAN_IN) & ((new_n571_ & ~REG2_REG_14__SCAN_IN) | ((new_n579_ | ~REG2_REG_13__SCAN_IN) & (new_n651_ | (new_n579_ & ~REG2_REG_13__SCAN_IN))))));
  assign new_n651_ = (~new_n313_ | ~REG2_REG_12__SCAN_IN) & (((~new_n309_ | ~REG2_REG_11__SCAN_IN) & (new_n305_ | ~REG2_REG_10__SCAN_IN) & (new_n636_ | (new_n305_ & ~REG2_REG_10__SCAN_IN))) | (~new_n313_ & ~REG2_REG_12__SCAN_IN) | (~new_n309_ & ~REG2_REG_11__SCAN_IN));
  assign new_n652_ = (~new_n597_ | (~new_n655_ & ~new_n653_ & ((~new_n650_ & new_n656_) | ~new_n642_ | (new_n650_ & ~new_n656_)))) & new_n654_ & (~new_n618_ | (~new_n653_ & ((~new_n650_ & new_n656_) | ~new_n642_ | (new_n650_ & ~new_n656_))));
  assign new_n653_ = ((~new_n580_ & ~REG1_REG_15__SCAN_IN) | ((~new_n580_ | ~REG1_REG_15__SCAN_IN) & (new_n569_ | (new_n571_ & ~REG1_REG_14__SCAN_IN))) | (new_n581_ & REG1_REG_16__SCAN_IN) | (~new_n581_ & ~REG1_REG_16__SCAN_IN)) & ~new_n258_ & (((new_n580_ | REG1_REG_15__SCAN_IN) & ((new_n580_ & REG1_REG_15__SCAN_IN) | (~new_n569_ & (~new_n571_ | REG1_REG_14__SCAN_IN)))) | (new_n581_ ^ REG1_REG_16__SCAN_IN));
  assign new_n654_ = (~new_n655_ | ~new_n618_) & (~new_n596_ | ~ADDR_REG_16__SCAN_IN) & (STATE_REG_SCAN_IN | ~REG3_REG_16__SCAN_IN);
  assign new_n655_ = new_n581_ & new_n257_;
  assign new_n656_ = new_n581_ ^ REG2_REG_16__SCAN_IN;
  assign new_n657_ = (new_n658_ | ~new_n537_) & (~new_n663_ | (new_n555_ & (~new_n662_ ^ new_n348_)));
  assign new_n658_ = ((new_n661_ & (new_n391_ | new_n393_) & (new_n532_ | (new_n391_ & new_n393_))) | new_n470_ | (~new_n661_ & ((~new_n391_ & ~new_n393_) | (~new_n532_ & (~new_n391_ | ~new_n393_))))) & new_n659_ & ((new_n404_ & ~new_n661_) | new_n538_ | (~new_n404_ & new_n661_));
  assign new_n659_ = ~new_n660_ & (new_n433_ | ~new_n499_) & (new_n391_ | ~new_n468_) & (~new_n437_ | ~new_n510_);
  assign new_n660_ = (~new_n437_ | (~new_n393_ & ~new_n395_ & ~new_n399_ & new_n490_ & ~new_n386_)) & new_n509_ & (new_n437_ | new_n393_ | new_n395_ | new_n399_ | ~new_n490_ | new_n386_);
  assign new_n661_ = ~new_n431_ ^ new_n437_;
  assign new_n662_ = ~new_n354_ ^ (~new_n355_ | (new_n334_ & (~new_n543_ | new_n361_)));
  assign new_n663_ = (new_n548_ | (new_n353_ & REG3_REG_18__SCAN_IN) | (~new_n353_ & ~REG3_REG_18__SCAN_IN)) & ~new_n664_ & (new_n349_ | ~new_n553_) & (STATE_REG_SCAN_IN | ~REG3_REG_18__SCAN_IN);
  assign new_n664_ = new_n552_ & ((~new_n336_ & new_n550_ & ~new_n257_) | (~new_n374_ & new_n550_ & new_n257_));
  assign new_n665_ = (new_n666_ | ~new_n668_) & ((new_n672_ & ((new_n380_ & new_n250_) | (~new_n377_ & new_n239_))) | ~new_n555_ | (~new_n672_ & (~new_n380_ | ~new_n250_) & (new_n377_ | ~new_n239_)));
  assign new_n666_ = (~new_n667_ | ((new_n433_ | ~new_n435_) & ((new_n433_ & ~new_n435_) | (new_n431_ & ~new_n437_) | (new_n404_ & (new_n431_ | ~new_n437_))))) & ~new_n538_ & (new_n667_ | (~new_n433_ & new_n435_) | ((~new_n433_ | new_n435_) & (~new_n431_ | new_n437_) & (~new_n404_ | (~new_n431_ & new_n437_))));
  assign new_n667_ = new_n495_ ^ (new_n351_ | ~DATAI_29_);
  assign new_n668_ = new_n669_ & ((new_n667_ & ((new_n433_ & new_n435_) | (~new_n439_ & (new_n433_ | new_n435_)))) | new_n470_ | (~new_n667_ & (~new_n433_ | ~new_n435_) & (new_n439_ | (~new_n433_ & ~new_n435_))));
  assign new_n669_ = ((~new_n351_ & DATAI_29_ & (~new_n489_ | (~new_n351_ & DATAI_28_))) | ~new_n509_ | ((new_n351_ | ~DATAI_29_) & new_n489_ & (new_n351_ | ~DATAI_28_))) & new_n670_ & (new_n433_ | ~new_n468_);
  assign new_n670_ = new_n537_ & (~new_n510_ | ~DATAI_29_ | (new_n257_ & ~new_n258_)) & (new_n671_ | ~new_n257_ | ~new_n469_ | (new_n258_ & B_REG_SCAN_IN));
  assign new_n671_ = (~REG1_REG_30__SCAN_IN | new_n252_ | new_n255_) & (~REG2_REG_30__SCAN_IN | ~new_n252_ | ~new_n255_) & (~REG0_REG_30__SCAN_IN | new_n252_ | ~new_n255_);
  assign new_n672_ = ~new_n376_ ^ (~new_n362_ | (~new_n235_ & new_n363_ & new_n387_));
  assign new_n673_ = new_n269_ ^ (((~new_n262_ | ~new_n437_) & (new_n431_ | ~new_n250_)) ^ ((~new_n431_ & new_n239_) | (new_n250_ & new_n437_)));
endmodule


